�� sr ,org.openadaptor.dataobjects.SimpleDataObjectj��d[�/_ L typet %Lorg/openadaptor/dataobjects/SDOType;xr .org.openadaptor.dataobjects.AbstractDataObject�]��� L valuest Ljava/util/Hashtable;xpsr java.util.Hashtable�%!J� F 
loadFactorI 	thresholdxp?@     #w   /   t GNTsr java.lang.Boolean� r�՜�� Z valuexp t MajorVersionsr java.lang.Integer⠤���8 I valuexr java.lang.Number������  xp   t CQsq ~  t SCHsq ~  t BVersiont 1.1t IServParam_FQNt >com.bas.shared.domain.configuration.elements.DomainVersionImplt PMinorVersionsq ~     t LBsq ~  t UPSsq ~  t Statesq ~    t VersionCommentst  t 
Containersur [B���T�  xp Yx��	|����ݕ�H>ۑl�q�;����@8b�vb�+�s ��G K�$'1J�)��R�BK������rߔr��B�Ж�P����=�ֲ��km���A�ޝy��?�{3;s�?,�h��<ڷŷh0.Z'�c������o����2��������?"�ɡX��P�_��`(v�ő�l��|1K��-��/Ի�}��J�˷�[���#��"x`Q����}gtAP�XسE�\Ñ�E�~9����+b-�Q��磋�����)�c8��z�hq�`��X��P���iQbX��a�*��ކ�.���"�E�R���E|�X2�7/=���ܶ[XZ[|�A9�L�g��x�/�9��Tb�WrR��0���7%sf�ƯD��d�þ�&(��2)�9"G7��=��^��6q�D%t(�c��ק䮰!��-�b���:O�o[s��\qR�-�P���8���f���{����݆��j��(GN���i���t+���b��f��������ִ�,��pߢ����f_D�Y���B���Ц@�`��C�DD���C1�Q9�MrV�ҍ�ͧ�+/z���,�aG �	�b�-�!�	[�HTII)���@O�R�����|+���.���6�'�R�㥫�<���Ej�u�7��c��Kt�r�eb���)�nd�.U�u��,o�'��RN�'��҂�S������4W��ˮ�c�����i���O���J�"�c'�g���J�<����1KA\iV��2��}*��įc[�R����\�U����!��u���]�}�Iɽ,z|1>�5�rdH/6�V>\l�5m	ҭ�5r���Ik��Jk}i��4�#}*�N����/�鴎2���?W���k:�rj�M)"NX�ԾU�G��t(͆��!=t$c��twj��KC{����}�^��<�%o�q7')7=��B�����z�Jo���m�	����8�tϦ�[��nIʭU)yZ�Un�L�Ӓ��*�v�B����֠�Z1�vH�,O��f^|a=FTٚC�=�qL�����=fO�4�����x�!���m1K�'�u���p(���J[�([i`Iv�&����� A V~�	A/� 8��!�Ap�B�����` V��Cp,}�Z� `P�@��`#G@�u���<:�ě���҂S����9&�k���Z���h�S�Y ��S*d �W�$uk:|���������������x���[��F�N������M��?�V�G��Y�����:�`�O�س^���C=Q^V���7ĩ��iL�դ�5�� oZ���z��ocw���鈄�\=)�4�ܓ<��:>{�F͝�76���E%��<�V����[�7�8&x:e���B\��4N���;��;BW�M���߻���Ѩ���RGI�@2ʆ����|u�Ū�b@n��G!���A�C�3��t���Vn��.�������}��=��o!�?n��~	�/ �)?��7��k!��� x�g!x�?@�OA�$?��jn��&~�u��� �!?��	W�B�)��3!�uQ���z�̕Z���:VTkT7�4e�NS��+T<�7$����=T{�U{���Y��ԑ���������;W֩n�B(vz[2U
MܫRC���<\o((���%Z�/+���]�9R?�4�0�⺿do��/�oT]S�H�}];��V�z��N� ߟ�o����T�v��Wކ�=ޅ�S>�G&A0�t�oB�����������kЭ[K��#>��b�  ���?���!�@���c�����k�	"� A\~��JI)�E�Q��֦��m���DN<�e�[L�z�T��T�tj �4��b�i�[5�6�uh���IaU����-u|�o�Ӽ����DF���a��,�C0�� X A%,�`wA�s!��+ٟD��jy6�"�X�j{MO�A���=횱|}ws�F�qz:�X��z�u�溓�����/oc�^���6�¡��ܫ��ǧ��0��h��f�������~ř�cx[��լ`֘��+5���ˏ����a���NcV�mkhd�]������
+���`@X�а�  ��
k+��`hXA+$�c0?��Ɍ?�����)v��|F��	K k�
OZ��*�AV�[��Y�-��rp��[�yD�ֺ�oWI��=y���x��(4C^�����
B������ޑ�������T�^���4[ӆC��V�R�;�d�>~�Q��]����|O)�RV<������5|������U�
�����	����)�����Vh���Bp'B�@IV`�z�Bp1A ���{��T,��`�z)�@p�C Ek�!�
VpXO�`߂�2E;%L;^9��������+:i�F��Nw�˭��튻�jҗ�Q��`+�
���zJ�V��?���������6��D�Iֲ1�	�![WꭺP/3?�P*ʫ��6E�ꡁD���&��3����uxe$��7p��0bk �����ݰ5�ۘ/��>�#�+�?&�f���x�
���7�)+؃V�ƬlX��,C+XrV����C�̶�B+XcV��`AZ�n���i��
6�,4+X�V�R�`�Z�����j{�
����2�������x��CY[l�-Yz�+3ꀵ�$:
�R;|=I����h��
Fb}����K�ܫX������1*����[���ڙ^v�1��X�X��c}[���d�ƥ+Я'8<X�%n]��Ҙ���8�`�/�A�G�C�?�`k�z @ #/�
�
Ya�h��
����L+8��h��S�
N+�EV0��Cp`uY�겂��
�+��V読`YZ!#�[! ׉u5�����Z�k���V�FZŏ�&�	Q��{�=�j�f����l�I91��/MBV� ��0Q���5��,����n��HU���$��]�ڕ���/0_��T@W �W �W��L {X`��W���!�p�J�W^�o��5���4:&EA{�DV{{�f�H��ҐOl�gӻQ퓭�A��mk�o�;\�W=Sܫ6��I�emT��%���Ǟ:�&�������Bֶ���ܵ�Шv�Cp���i-� ��j��N�f(�_@����Lf@�0�[��H�
&@c$���TC R	`r`r� X
�Wx!�� �����I���5�5�\C M� ͒ � � �� ��P� 0��=�i��!�$�2_L�Y&��h�C8e��^��w�����W}s���0��	�tm8�hV�C  Nh�H\���I�I` -@����6h�;|!9�*��*6L��Vc���ƞȼE�.�pE�63�r(�
��n�ӂ(�әc]�J����k<�~���T�;���8M�駦f�I	��i/դu�|��Ѥ1N�iYx��Q���y5���&
c��B 	0j`6K �J`u)L/�"(� �� Nf�
`�	'@Ղ�">�H�>����J g� �� �����`�\'��^�m�S[g{�!��l���[��Y��l&��_ﳗ�) �G]њ�@�Ǒ�wm+��׬�u�t����nn�!~��
�-O�c�z�
Vz��5�JvO�d���L��Lb	0�%��*�D� #J�j,ɕ��` ���w�/�$!#�x�6A�{9߆�{0P�� �#8J��@ V�p=�n�B���=,�Jޠ�8u�g]�c'�wMAJ��m|3 wVi��m�>S�'a��tlH�w(� �� �� � �� � � 6� ӓLm
0�)��*��*�|)�r4p����~h�uj��j�����`^~����=Y�#x�0�0�0�c��
o�#�
'u���uz�zzqAhԝ��{S�}V���G |��v:Q��~	_`JJ�))kk�eX7��4�4�P�f��Ӡ��i]Tl,�� ֧ ֧ 3s��	`�ZV��&����Ѡ�/`Pf�{�kf*:4�֎VUfӷdL�0�(�|� ��R
�@E`&R$ܿ��	ʪ�f�/�»T���N�!��X�����GG��頞��z:�,J��;bs+�NL\��gHʍ��;��К��K�5^o�J���f�ͪ��.~vY��ӭY��ml�,$�rm�H��J��n��`�X.������U8�A[.RVX����u-��P�_�O�a�Z���o��-/@�<�5�� I
����-B��l���lR�[��n�^��z)f{���0g.�KxD ���,RX�!���5a:��������	@�/��/��/�+@�iQ��+K��|��$E6������^��/�J��:�)�"h?VϠ�@,��A��v:.���s`� �N�"j"j"5"����*�Q!0u��D��2��{˷�&�s��_E��D�x����r0ga�9��Ȗp
����!��yX�0[O��?��0=��àf��뮙�̐��v��[X�0�-`����m3�f����h`]���f���Cc����&�9�����i�H��!(��]ҹ��5�I6M�[�<߱NX�#2�+H6��ʴ�M+&,�I������}��<����vX ��q��%#B��P�"�(���P�>0}Z�"C��I��z�mܟ��]=���\g�"@(6B��� `�A��Jb���6g*�g!�Rb[R��Xz:���Ҍ
�ꍫy�;SVq5�^7�z�U�"�
a�D�iN�5"����!B�&���x���tF�����?#;P����>j��ԡ��A�X�r�nt"�.�.�].at�=����Wj�׳,#E��m� ��M�j3�]�[2�)B��!0]@ M�n1�a�E�A�돰�-��I�*S��]�F�^C�I�m�<_-�WZZO� ZI{@ܝS���^I;=��J>�,Z���{��nO�-iU8r,W;
��Z:V!l���b\syYr@z�����,�SP�,����PץK�N�.�|�Q����$��x-�� ��������r$v�xw�m]�TF㖮@�n7���	��@p��P�j���-�Mx&�E00DX�,�
]Q#|O��9�h2w4���X�U�"�Ua���DX�,�E��&ry]���C�x��t�+f�����]	�^��h�:��D�x/�#ޏ��@����IJkê��I���;�T�m�L��ڰ��Y�[���|@���0� ���sŧ1�)��4;,�BÖ�	o=N�7��q��VBL�G�f�C��U��vA\"8>Dp<�0%-���۫JV]�U�1��5�%�*Z�'��r$S���0�?�&.�)%�7�%�y5`�8Bge�w���#z�4�no#��ś��Ya`$�`$�0�,¼�˰Ep�`q�0� �� LEn�+:�H�HAW}|啶�I_aс�>�f�R}�[)�z�[�~�-���Ґw[��
�t�K`cK0z��4��k �.s+9[R�^z�Fr~����2�e �B/������\ܹ"8�Ep ���q'%<��E0W�s"sU��C'�&�&����q0�Ef��~�-*#����I���Y�6��2�e �?Ed�f`� ��.�sC���"�O� B	�",���#Z}�!f�$L�0k,¬q�$c�� 
��TQ��,��`+ici���{EϚKE�/a�L��2֕�0-�hJ��w|��&���Y ��5Q0&���{�Yɥ�t����������u��E����Y�a�^��v��E�Ʒ0u,B�X`��R��{��G�v�m=L��c󕸧�~W�pR�Zl�ʹ�Z|E��<������t%ФlK�P�R�v�$�%�HXo]�x��r@gR2&�`Ĳ��t_�'wyX���_������=)��Y���b6���)E{F���h���3V���/;�s�Cшerro��'俯������+X����X��1�:Diwk�2�����ɻ����9�{�H��W^����U�i�h@'H^��8W�Ep "!�'۸?�`�D�`�,NH�Ek��K@g�po��JK��MH�u������+�A������+uԭlL�_�2>_W}|	$I����Hɉ]�ɿ�Ǖ?R�鑘�Am\����xt�tW&����2�
�i]�\�����`�_M���V���N09��v����w
Z[�M1խD�Z}l�xG��Z��1�H����'��m�`8*'� �|����{\�Gz�	�-��mz�������KWu��t���c�Ԟ48\��Ba��Ӹ��zM�@b𠚆��#4�1�u7��䫿?����y�R�Ԝ��U�Uwc��{Q�:��6���d�D�`$&}&��뼰�
�0�H4�s���U�>�P�K�R]y%u����E�����������E�|�?�v����T�q��:�k1C���`0)�`R��ҏ�ؤ0M	�|� 1��$���`�(]�
�`�n	V�H�t��� �%K����!� ��*�k55�_�ox4�c4�[4�>�u��گ���r�Ǫ��4��"im�n!�ʢ�xB��L�J0p�`�.��rI�D���t�+�ME�ƶ�H���$p&��/��ړ��$�
�-�1	�O̻I0ؖ`�-�҅�'��)�ר 	��hH`kH0I'���`
k�$�N$�q��C�H���5@�d	��,,M�XN��PS;|��cHLv���In������wj�x�Wv�&\o�PK�� ��\�őPP�ok[�}��\?����Wi[��BL	>Z����Iz�yH`�I�a���(��
 =�IK��J�d��6b�R�R�b{�H��]�oH=v��K]�t�Km������}+��X�Iv5�U�|�-�%��-t���>�_�!�W5�x5�/��a��ã�u�/`-���zV�0�d�9*1S̑��"�� ��"�m�g����6;�l1u���fC	l1m�$�)��&D����=��a��9*^����
�/��U�T��N�B�
3e�0�^H�w��pf�$k��c#��F�Kһ$�_��Ho�Xo���B����H����$>��$��Az���S�Y��r��ч5]�d�Z�^̛l<T�Ki,�XB$�J�[�ۗl�������K];�1��z[j�0p���lp���,�߶|�A���?�H����!yp����pl�~ u�A,V�t�=��2�r��_�����2*��FpJ��lQ�����_�8���������.�w������-݁P4��e&Z�F�r�>{�&e<��_P���'�������~�������)�S)g��7�_,�����!�+�0��g^RF�L�Z�d�s`I��:)���/#�\�2����hV�@�lცQ\��~Os���	�[��4T�l�f�q��_�*z4��+7�Pd�2����������mM�)�����ڵI�I�
T��\�`6�V�*��ʷ�j��
�-GU�@%���%�[�� ͱq$����ioI 
�z�-)H�EjmV{�tqI��p �ĕ��\�_��i�5ߚu5���@�غ4����X�ZZ��fj߇x�M/�v�7��h�YA�/���z/���J�����B���}N��t���a,���F��0ڊ��@M6hIXO�"���eS�-����+]l ��t�>�6��ێK���E�X�Z�%vC��Zsۺ��V�-r6X	e�N�V�,4���F�� ����Z��hہ\���a�ҶY�m"Jz�'����zZ[7�h�#ض#ayC]?���u07o��ð^^֨�O��X.�˃T�ΊD�g��k�\ɏ`�Uɬ��k�0�|������
���E�Ì��3���pg����aU$)��S��K�{]���fm�Q�� �1G'�O��g����ϰ)�Fh{_���d��k�e���=����Kb>��=HYy3m{ �a�k�Uf��o��r��?6��?��������h�l�T/F8�m�t	˕m[TO&g���f�>�ڎ_�����&�'��&��U}(��Hժ_���j���~ߘx�U�s��n�Ŵꈙ0F�`O�t�^�'��y����-��=�����3�5��b�������2*��Fٌ����/X2x#�3��;����k�j�6Em�A��}s�P%(r�͢�6�L�<Q�4�B��b�B71Q�D�6�N��5����¸>㧢�:t�9�	�}�[��d��|���>�*'�	��AW�L���5I]Nȏ,O��r!�r���q���#ד��u�Q�q���G��:�v�\'���]���#ӎa�t��c&Y6�5��(��y�'"�byk
�\��+�b�Po����IPV������_F���(4\��:�-J�����<x8ǚ�(+����,�QgYB�A�_�e'.�=��rw?��q�V��v��v#�A�6�wO���!wB[�P,K�f�7L�Q�GG�����i��R��X7�`!��žW*D"Z��lx��t�_̲ߌ`�2�#k��u���hr
B�J��x����)�����}95b~�7?��Q@ܚa�nNs?1]�h|��:Yw&�^Kg��*�E��w ��PB���=Bv�B����#ە�fۣ��zs�(�?m~d�j�Z���Y���^9���0>�Su�_ʲ��N�-�5���@��&�5��ɕ�2���W�45Ldjh	��2�έ����P4�2r�������=A�ɯ7�f�0���u�.��=vL!�:�^����Z��50&�L\����0CG	.��rnd��r^��C#3u429��1���`�C����Y:jp�ԐKؓ
ȏ����|�q��m�ړfxk�
�訠0������`y�����:�Ot0�Vۓ�)�?�ݝv��x-���Bib����B����@�ŞG-�|ML�k"��܉,V%ұ�x���z���y=��MG�"&�Xn��q�#�`��@�b���uoY��s��p�쮣�b��1�������[㵲PG+���;o�����y�����>
㔰�9�
���j��Eöc1�+d�O3�3^��0f=ěW ,�����a_i,�E7�#�����R�f`���v�Ax��^�r���g�N�'zc�P�/ғ&�c0���f�ʞ:B��䭵�}3{�؈=qx��ҭq�ؿ9!y�.g�EOSI���H�$�a�?����I>ax��ё|RC�?ȶ�W����k:R4���	�*r��"�'r�q�`x��ӫ���_!#/*�mx����Y���X#�..{���\G�r�f_�W��{��9��7S���:(�Ecr_mt�c/{���GN�뽃����~����Wc��-�e9ޢ;��`�'�
�)�5q���I�f|�BG����h ��0��~�_�m���@:��(>u:�(����|V2��+�&e�g�^'�0��¸�|�xtr�ր�.^�ǷҴ>:y(��D7���*���eoԑ��%������=�^������w���(�����(����_��C%�Wav�-�({3&i_������v/fȾ�b��L�;P�vT�}5��ކʷ�h��(���P�9~g�]C�𮍡�vc�]�_����0B����{�$���]�Ũ(������y�%(��;�!��1+��1��o�:엡b���엢���L�����hc(�䙶�KdfW���<b�ǚ6��5�]�߻��7��o�������av�/����c��71���QL��1C��0+��1��?�:쯢b�/��쯠��/�L�Ǫ���oW������o��1B�B|ձ����:f��30I��y�ӱ;fȱ ���3혏�p�C�:f��sQ���;���٢�������s\��@�qv��e��W�#t⫎��$G ���CE9��$[0���a�̊#��v�:��XGU����h@��4fY��y�1˄�([���N�����ւ�p�A8�V{��.|)�BVN���B����m1K���Y��_�?�]9�I�JyHR�0���,�i?�8y��@�C�'ů�J��Te�ɚ��q���ԇ�RZ��к��ZRjIyh}�C������kX�����N��Фwsm3;k��Y�N�^K꽉��PH���TZ��Q�Р����JsSZ۬�3�)��F��r��&졹�M�ΚA9�Xu�=,.�o�knAL�TP�y+��콫�A#�(F�x_u��Jr���x�x�t���w<�b:��9�Ŭ8���v<��p<��u<�*s<��w�Aw�tmVZh>�V�KU����kk��cQ�ڈk�Z9X������dpl�!�ԑ�����e%+�nK|E9k>0��Up��� ;�`T��Y�of���t� ��P	p�8���q��".D�p��p�Q8���01��v�_�.8���v�韎�!x�����a���u�/��ǯ ��B�)r0G�og�8F�qWB g~:~�*w0q�Q�������sfpά�Hp��)�3ep��N�e�Nu�)t8�.��G���:n� \��N�q>q��:�U�`�|h��(SX�ꀃX7逳p��Ku�����a���dA�d�y|`˾g�4R�U��ҿ�c����ѐ�7����m+���t�2�T��:�H��ż���őr�㓁Ò�4��(���e
�)W�<����C�6᫅�PI��cvBE.�$Wb�F11C��Jaf���QX��-<UV��_x��x����j��W�?ˮ��r������W�G%���-<Ux2&Yxf��t���P�Y��³1Ӆ�Du���-<UVx*��i���|4XB<��hS�f��|4%�tp:������c�@ܖ�ĵ���i>(M=w�=t\�M�i�^ �q7͗��gf���q7�'��gR��'���i>M=�	�=g\�M�h�M ���*n��CS[q�Wq�|�zJ�{۸�;uxqS�7q�Wqk�7�P"��q7�WV���/���i��L=��}{\�M3"K=@��h\�M��f�4J`2�dl�-^��3^@ܒq7�G��'�����*n���LW��*n�O.S�Oq��L�,�%���e�;Z����n�W�~�J*��[�STT�u�d�m����Q̢[0CE7aV�n�L݈�(�[�TY��P�E?����e��y��y`W�7��߻a���jї����0�E�BE��I}��/��,�3T�	f��S�t�Ǩ���b�>@�}��/���-w5�;�k�v}od|�W�FX��W�QI�_��/GE�I7`�@1��1C�+0+�u���Q��b��G���/�o�疻��]�߮�o`���0�����sPI�������*>�,>3_|
�Y�M�P����31�ŧ�:�OC���*+>�_�c������>����������1�����gPI�`v�AE?�I?��/~�,~3T�8f��	�t�Pŏ�b�F���_���ǖ�|��PQ�8.�}��_3~�>%9��g��=]�$�$F�f��\�x/ysp¹�?��0��W���0��W0��?m�Y\��T��(�)�,���@|S��x+�U�K7f90��Zё8Ld*)�L�yG9��ƺ�}_�K����k�Obۓ÷8O�ٰ���dnY֙c�6�,���j�ZZj���p_���x�tmW�����FoW��ZxauZ�g1�[�'x[NKB-���=;y�ry�X�����3T��U��P���ߗ&S�����ȅ}T�,Q�����B�{6u���TQ�p�a/�[�T�T��_���>J�W�XU�"5��ѧ/���ҿ��<'�N�,��K��ݣv���kÛj�/;:��࿩Ҹ�w+T��*q�W�zj�7�gia��R�?ݲ,��ӭ���R�,����V�Q~�UÎ�I7�������	l
�=ݱ@��ˬ�w����Z��u�W9y�Um{gCcgm��ꛋz|1�{���S�����λ�sΫ3�;=���*K�^������+N����z�z��vU�U �mt�^�̯j2�	;�*W��܌+I�����TW���]dW�
�[�5Q�7[K��WJ���J�h�Q��N�p2�a$�+#����	{5�:��IW��I��bC�8�1Zӷ����G묍�_ϴ�����#�q��lG���J���P��60�-�N�w0苀D�U��!��س%/+e:E�Ÿ�]C�r�`!g�b�]���^x���u���v����k0
mgl�/V���j}~8%��n�R��ͭ����7�6�/��Vi�e%j	�!�HL�T��yPTDi< �d���*�.��?�4�DV�^L��������K%(e='m���Gђ�C-�GԒ��Z�(�LK+IR]���4��c%��,y!y���J�9	_r�YW��N�S�W���W��E紱d>N&�6�d��9�H����`��|���W
U�4+��̕ZFJ-Pu;�Ԫ��N��m��+�iT~Um���uO>�E���0'����}_>��yff�x]�S�F2��U�1ˤ�H8&���}r�
{:vu���\+G�4ț���{:W}�(�>k~uQzoN��V�}��G�x< ���A	���+X�س�V����R��B(��S��4���v��7:����5���Y)p�C��	�0��<dة?h��p���^�bq1N�hƹ��s����D��0'��d���KNؐ�y8�)���)b���2oRWP�Z��>}xs6�p.�F�(j��F� E�02$�V���X8�d^����O��2����`�Q�D��f��PoP��G�	Ï7
z�b���lp��R`�`L��=6ц�ȪI�8L��ʨѝ��Nu6�\
΅���ܳ-���4�<���SihI���(�a�T:"VA��t�v5����.�%_��Q6I�C���\3ߑhZ��6��Ջ�^E�Lڅm)AJu?b����+���6�3����q#_L4b#���y�6ƌj:S�w ��֝�VjY�Fz�)<{/7k�TMkS8��i�9U�`�����lI��X���VW��m>^6M�=Qy�f����Ix�M#�BU
p��jB��L�{1%ߞ��@����z2'�,�����I�u�SS�Z�������"�rs�&7C}����m=��O�h�3ɜ���������okj�ޒW77pw�j�����(H���S���ʝ5�Q�Õ�r���s���	��:a��-N���	���)`���	��J�B���?Q0͡M��b뚛3����:^�q5f�:aSX'�'�V)�����5�8�GO@x�\�^4�$��3�,�o�N:��F��=��N�����T�	�*:�#F'l�ꄍ^�-l��
�+�)'lS�um�����u�f�lٔvlu���N�t�	��:�Ŝ8���ivޅ��	�=:ae��~�N��5DN؇�	����0�	�M:o�:�k�|�NX1��WN���	[�:�J'|��$'lX����N� ���hJ4-l�Xv�`v��������;0v�V�r�����Y��I����Î(�A-�YA�^ڡG���˧�p�ߧ��p�L�&7jt��_���?S?��PMr�!>�1@M���4Y��4}Ÿ�IjP�d�����F��%˸�ȶ�8�BY�4�WR��*)�e|WF3ӹP������%�o�;԰�%��:�j܄�PO�/�J�Q��X�&h�I�W��P�U�y�ں��g��/�����brĠ���Y��^q�;<�в{�f���y�W��*c���hi��4r[uI.�`�Hj5�=��BG�敎:��2ct͢����h�[$EGK��Q$=�O:��_/�����,*���T�جm8�e��3|w�f�Xa�RZ_���llj�ll�4vw��f�.�h�l�ʒAY���3&�����}a�u.��F�%s�-�yP��uc^�,�ӭ���,�u���@(��vd)єlN�%��ޘ�V6&ġFzc����ūi�=���j��cSjj��4����c�8k~+*j�|�\T;�f�̥�
���~c�"�F��}�TK�Y�7z-mˢ��ki|[��C4���ҹ�����R�נ����j�U��ҫ1�ҫ0�����IB�l����� ����X%9��R�ҟ�K����R�қ��~E�t#��ڥް#��v�ZA#{KU �񛟺Q,�bQ����K�,Ï��"�<9Q]c��1Q��ay�:�����[(1S�=�R�ǫzP��D�J���/�lM�K�v%AO]�Y�x<@:���J	J��_��7OV-�k���X��\�
^�T>MYg�}�:��6�|oyI�xA�o(<��>DX+*oꈄ�3�'�3��V]x�'�X`����&F
-�M����Z���5��^ANt�B�fK
-��|{e��_ɵ`���k�)��2�!nr-X�W���5�_��e��Z௭5����Bl�0k��=>�|e�1ڲ)���"L��)s��e���27�����2'���3TV�Y/�_^�Yb_^ "r�xH�� �u��<�Ԙ@�==�JI�5g��u��S���.t:��ٜҕ:�R�k�j���Hb/�7lu�-�g�����4���T��2p%���\�'p�v��&�ʖ@ g���ڭ2X�U�����U�L��@��
W@���I��5��%���U��VS66������Z|堦�1x��#+�.�5�ny4��羚:����5��$;�^v>\v	����ӂ2���5`��`��2�U�,��meM(BY3�l���IJZ���<�Ŷ���y�m��NȦ
י�h���͢'c<�6���b�P_/�\k>�d�F}�Ls�W�u�Ou���h7��#��n�:z�Q�D���2Ҍ��oJ<<yݨ�k+Ǩ�����T��$� ս>�{a,Bu/Fu/��ޒqE���ǀ��'���ӈ�Ӊ����D��D��D�)�!��?����q)�r1>!	v	A�/����?!�D�_M�_G�_C�_k�2��[��ߐ� �o'Q~I��J�����k"��|!~���?J�������������4��k<�����/�(/���ϑ`/�/����4%�����'��FĿKĿC���4Ŀe<����V�"�+�K"�S"�s�?(B����,O��<Ōė����e(Iy1�X^���OF��KP�r�Y�/W�� ������$�tL�|&�R^��*�F��kP��D�,�l��|!�eS�7����_B��E�/#��4�{O<�I�W��D|#�!��OZN~��"���_�/��3%���C��."�Kį'����LC|�������I���L�o"�7�=D|/ ��yB�3fJ����[��-D��D�6"~�4�G�'�"��"�,"�L"�T"�t"��D��D�iyB��kMI��������&�K�����4�_j<���7�?%�o �'�#�B��������q��)��������-�D��D���;LC����0�����"�"��D��D��D���B�#�$�"�M"�OD��D����׈��MC�K��"��$�?������w���������񷛑�)��)Q�)"�8E�Ԧ�\S$�h��4�e8�S���JcJ9&0ō�L����2şR��Mq�S*0�SJ��ҽLI�nD��D�\"~����G��7�SfO��D�$�׈����}�����}������D���B���$���o#⛉�UD|��4�7O�:"���8��?��?��_O�J���?��ߐ'�O^mJ����">H�Cć��>">d�7O��q<",�"~�=O�/�`J�/"�/&��#��%�/$��'�/0�gO�D��H�+���W��%�O��������^��)���K"�"�f"��D��D�m�!�㉿���ĸ��������������������+_�?ڔ�?OĿ@�?C�?M�?G�?K���4�?a<��'1�B�������3�&�6�7"��<!~��$�"�K"�"�c"�s"�S"�3����Ļl����pM�\�(�ˎ�r����(�ˁ"��0��	�B�{f$�5�wբ$.��U���jP.W5J�f�]n㉟O�/%1��=��D��D�""~	���x]e�9+lQ)��Y�zxa�'l���k��ڸ�2c-j��]�(�k��Z���V�\�f��u�����Ī�X��\k��vbu�ZO�v���j�n���ى#���b2�_�.}�~��k-�b�|h�\˷�,�S�8H&�@_�����T����h�A8�ޤ��T����o�n�rh���������U,��������,e�ܓ����Ty��"&���2\��D����SC 5��H{���Z81]�h���邅�.pg������h,���� c[��5�:a-Al�ZPK5�&9T��HԪk#A��p���k|]G�4.�J��y]2�G�؉��R�Ay\� Yr_�j#��z����I�:<�-<��n��u����]ے�Ym��:	_q����vP�'kvL�?ڴ��9�?���Llm�J�, ���c�Jlj��
����Uv��X�7F�T����ƣ����h��Puu$/��ό_�e���Tt�����\�^����8O�hjC��+��C�}	�:^��g�	����1qB�0�~Ȓ9M',\Vu������5?Ku��������n�}�{�e��܁�ے'���W��`M
ɉE]�O�Y���B�ZZ��^��~Ou�^�{@�4��|� �c]���N=�G�N[�C�RZ�M��I����D՜�P׶�[�Tح�CR�[�*��#�Vg�F��Q�`�tO͈�r9mm���c��EO�&�F>��f���Y��r%��qXʭ��hܭ/����dN a��vp��.�y�! �/�`}�֜�G�������eCLָ����F��s��<��\�Bs�zU�c�C8�\�q���S�RU�fu�"X�h�/��bx.]�=s�� x�]�pv�z?,tA�q���������B.X��zK�;x�\���_����Gt�i�%P�����
�L�՛,xY�%	�I5�*}��)`���]����~]s�*-��A�L�5���q)t6��kR|J�����0���Oh���v����D�����g�k�n��1�6M�ٯ̎����)w����+<�Ȱ-d�Mf��Ox%K�"�~��+ԋ���>8�?��{�3��64q}5�.�2p�:C֯�`i>�{]?�vbٹK��$�]�4���X]_`�K�,�Dd��at�k5>$�R7KÊ캙�I{Ÿ��׍ȕ���RV7a��I�;�7[�*<|X��v2`���7�xVI���u;��.B*ݰ���I7�zA�삏ظ�_�����r0����d�gi?\��`�=KI�ZoK�6ܵ��w�W�11��vw%C�z!#�A���ܱ�,��]mE���c;^�Ð�+�%7��8���Hٗ�r*1���Tb@2���$�����L�l��B���\Ͻ��j��H����+�b�Po�M�F�"�63j����K�.
$�� ��TG#ksV��$c9s�b��-�� ��o�n��X�$�P%�M8f�� o�lF?���%�Bx}�Z�D��2»w�p �E�od�l�#���g�|����V���D���˜�Wc��8Dj 5FY2�t�)y-O0��@���!�0:"�O$��A���oK�c�d��'Uu\�T�1KA�jO8c��$�t�]��W�*�J;Tﻕ�&b_�r��μ.�Ơ�I�_C}#w����g�iğ^-q1LP�Q~�7S�6�fg��N�o��=#6�npo�au�����ϓݰѤ���3p7,t_���F�.e�#zC�����P���z�nu�ުK�ՕQ�C���|9�{�8(��7,�s�������zt�8=���M3鯀��0+��n؇�ͬ#���w�n��L܍T�`ҏ��ܰ�k���aq�2@7X�`��aZ����z�vn�*��>&w���_�ѥ&��4��X�>3�f]�����V�l7nN��qÄX	x[���X��ɑrR����ڙ\w��qc�^�ycx�t�"V+�:[gi�=���H��p���+�LUr����.-��L��@D�l�x�}���и2l��ً�G=���_Ƽ����Y�8
k����?���>�*��މ4vVC�8_%^�!UY&b:�ʒy���dĩ������dx���c|f��ᚅa�����a;��k�r��4���μ�*�\)Y?�R�}���`�{c4��)�L$��㨡��^����b�7�f�?���Uθ�qszڇ���f���&����c�BQ�8E�]�c�����T|_�8�8��8B�����H��'����!+��P��!��$��$z�$Zo����K�*�DL2�Vz'K-���#���:�~0Y�JNV��GU�SUbՑ��'T�<�zLu�#���䟴�$����(}!���0G��˪�^Uŧ9������7�.�����r\� z�� ��]�����~��ڗ��_%��ZT~�	�?�I���Ƶ�R���INǈJ���	�_���D�m�|��Q���PƊ1��[Q���Q��[���D���k�֢W����ĸ��E��3U�;��N����>�l���)���#���$�,�4��i���������+����&��g"�/D��D��yB|�lS��9�o��GD��D��D�'�!�É����B�r&PiGQ*'b�*%�� ���"T:0���|!^�ß��WN��+kP��J���S��F�*�P�ʩf!�r����%����{����D�B"~??_�_eJ�W�uD�D�r"�`"�@"� �����7�$F+�Aķ��-D|;���_�/��b�O'[W��t�u%�l]I'[WEě�d�J�O�����+I:ٺ2J���֕t�u%�l]!��d�ʔ���:�=�V�ۑ}��hg9|�@�<V��_n�[��Y�+i1\�I�X%-��ܡ�|.s�;�3�غ�R�>G��(��S)
�.�.�_��_/ID�D�l�V�W��]���9{�es	��eT6S��jz���,�]ڶ��&0�w�~��N-�a��#[~�&�j�O��R�9Z�S�c��f��:��'��~7�b���([Т���1�f��������"���1�d1��o�" [��,�����=�=J��N~�Yץ�`3�i�s+��(��7{(��ܫb�����==���jW�ڿz�<Y(T�4�̨
Dc��r���b�B��|�����2���|"3��#a���v��\�1z�e���^g�Ng�[��Z���#�}��|��-�W����v��������{me�F�jrN*f6��x ��33���j�R5����V����2JG�-�!�Q��d���r�L���}s�r�j���T*K�T����3J]l�����W��,�D4��g�^�Q��R��ٵ�F�J.��LQ)�;$+�1�C�j>_uJRu<�Xu�Vu"�UuJT��8$����9$���W]Db��	T]��T����:ů:�:E��3[uv���+�cJ�&�D�_I����!����������q3+�s"��|!�S� � 7?/�i���x�'�'1�&��H�?C�?A�?E�?K�?G�?�/�?oJ��F������&�W"�-"�m������������������������7�)�9�Q�_5ٌ�O-���$S'��S'bjSQ��v�h��,�O�N�T><u:�Q�	L���L�LMu��S+Q���(����Ԋ4�l�>�XnP�f��L�3���&ϭ��g6uw|e�����(څ9Yn����y�a��]�0u�і\�mO7uE[���h��]{��ƴ����/M=<G���%� ��uY�A2Z�4�����$a*K�������Xc$�8�e��cY|B��0b�c���ʦ�r���:k oVL=��=atۑ4�AÊ+�Eq���ₘ��\^�ر������P��8?�%��{�Q��v��6k,�e2t�ힵ��m]�]�v@�鼜b�� ��zU/��d�R��P��]����:���r�P�U��iI���甅�f^�#֨krQ�rU�&�Gz�����&˺�ݐ_�D��{��L>�wU��e~1���$o���=�Y����Y����ꢼRT����˽������$�~�Ee�V�zi>)�������k)���<����%{S �n6���e��PkyM�oU�_�-�f{�U#�^ս��UV�W����&��rsUo�W���Ī��h��۵O��ۦ�l|������>�J�<*�Ө$�صO��]�ԍ�8���NQ)�O�WO7�|�S�|��(I�(O�aj�O�\Տ�D�O�eR����A���/���o������T����~ů~�~E�~3[�J�,C�^jJ��M�L�@y�'��/"�C������O��bL1�i(�4	35͂�OP�i6a���4k�_dF�U��ӪP�iSP�i�ڴ
�k�%��6��&N���D��$�\"~?���E��!��������$� "�@"~_"�kD�r"~?"~�����7�m$F3�B�B�7���D|+�2O��z�)��&�"�'�#�$�N�a��O�f"~���a"������!"���?:_�єğDğLğ@�O�� �Ağh�5������I����������s�������s���)��%5�"���!����K�"��D��D��D��D�mD�/������LI��D�CD��D�=D�D�}D���!�N�����x�����������#�<�T�_�kJ��NĿCĿE������6�W��g�����������������������������w�?�b3_S��ה�$5v��f�VS�r�8P��B�_S`8�5n|���ĠjjP��j�TM�_S���LCj�cfk*��j�)�_J�/#�� ��K��ED�b���x��'�=$�AD|0���?��_A�����z���kV��'�5���.մ�+5�XM+E۞�O��z���#�����F[6~*ZWT�����鏚�rw$�3菱w��N~�\C��֜����k�'[	�!ݏ�G�i��}�5�'�l�rNwZ��JV���+zW��[C���g�A�s�Ù�\�b����̹�n�/�m����0dK��k�"[6�"�������g�5gs��#"�#=r��=4Hs�g���y͕��\�Lgk}��B\w�o[�o���}�'�7����7�/2�!s�9�d_l0"���H̽���)U�;�]���~����@NC�M�쏚�sĜ��ʥ�����)���^���	�.��q�%P��RCN��>%?�U�*�|ݫ塭Jkd'g��y���ʦ�6�rz��X�ws��?�U��b����B�#�p?^��n�Y��,ɥ��p$�,��Z?jm�1���i-�c����9G���">�1
vƨ��,�l7��|�T�ͯ�9���;D'�K���4(��',X/z7ǌ��V�WM��9����嶑s���j�WgdAۥ���u����bc��Ҳ8�j�u���d�4k.U%�����YY���<W����A���S�n���0l�b���Fݍl�N��]���6Ǻ�_c��9R[�Ǻ��V�^�}��Z�`��A���۱�;9�]��j���Ac�7���jmy�?{�u���`��v��F�j+x���d��m�o�2V�u
'f��ny�Y�*��!T�ȝA�9R�X��rL1F�t�6�h�#G��y7Zǉw'�7Fo��Fޮ�֟#�9���L�φ=_:Ӯp�gPgz�0�FnK�t��F�$91p�Bog��&*C��/d�z�-��� W�
������Fv�se�9�,��D��#�*�����gw�:�4O8+�ʾ���sGg���򴂲��@�\�Y���9����l�=���hkj+���ikL,��(�@��72�l�#/9s���O흂��Q�Q�+._5�k�ߠ��P����䧶�f�`�qf��������9��cj����ǹ����Ì��;>�\[��oTOzl
ۜ#��AOZZuw�b�������ˠ?ݞ#��?MYA����,ԧ��$O��.4Ed�����Pqt�W�˗9�It��������`���Yr7��ɭ�YT�]����(·+���:�;�<�:ĉi�0䌫R�
��<����ȍG�sxNL��JҘ#��y�$N����o�b��/b�	�/vY���T�h/�(�䵘����j���F�<2t�P������#�����%{�fv/R��A�D��[�!F���0���=�K6�b'��x��	�|��|�RսXdP��2��:�ci��0ga<A���Twt������/9�v���K��#Ʒ/;~�K�7��G�)�,Z?��V�u�/����ci���%~��Y2Bjdo�)��u�h`cv�=�~�2�ys6�3�93`ܒ������������L'&6���Y���aG1KqcGD�*���8����G3k�3@]98�h&�2s�J�J5Kf�>�3͛>ui$b�;�(f�Z}p���G1K+���֔���ߓ��}׾�J�j��t���~���s͸O��c���A�df/�8s�6�h�k�f�hf�,�t��'�ڧkf�y<����E�9��bU��?s+
6�Xa�q�ٙ[�dg��SLI��D�yD�7��3��s������MC�i�%��"�{D�D����ˉ����'⿝'��XbJ�o&�o!�F�_O��D��@��h�l<�&��!1~G��E��A�����-'7�yB|͵�$�i"�"�q"�D�SD�D���!�Q��������:�
�'"��D��D��yB���LI��D�'D������������'~��5	Ř%a�&�(�l��YV����*@fM�����ڧ�H��*|~I2˅2Κ��ͪD�f�Q�Yf!~V����"����݈��D�l"~.���ߝ���'�O0%�����������MC����Dķ���D�j"~%�Lķ�mD��|!�US�#�N�N�w�G�G���� �#$F�Oć����� &���c���<�w��D�)D�7����������!~��ğM�_Bb�O�_D�_@ğCğG�_H�_Lğ�'��v���k��k���W�?"�H�_m�g<�7�"1n%�A��F��D��B�����%s��)�����������������4��e<�O�/�����$�"�!�#�_ ��⧷���w���o�o�'��J���4Ŀa<���!1>%� �?#��M�B�N�I��'���̌��.��g;Q���q�S�]�r�.D�f����'~v><{�Q�	̞��̞���]���&�fנ�k1������WLI�2"~O"~����_L�/1�O�r"���8���'�W���uD���?0O��.����D�:"~�A�w�D��4ķO��D|/������x?�M����"~T�_{�)��F��1">J�o%���-�!>�q�a�� �Ib�JğAğFğDğBğNğIğ�/��LI�w��+��ˈ�K��ˉ�o��6�O��D��H�����?&�D�_K��������&_����������5;�["�7D�����_O�D��$�#D�cD��D��D��D���?��	��O6%���/�/�"�_!�_5��O�߈�����$��#��N���������'O���Č�ϑ��96�d����
S�#�\s�(��4�a8�s���9.c�dL`N9�2�35�ş�D�攡s�`f������yD�|"~�8g&?���M��1�s�O�"~?c/"�kD��D�R"~O"~"~_"~Y�?c�)�?��_M�7�D|3���_e��'�K���XO�F�o ⻈�uD��D��D��<!~�~�$����"~3$�&�1���o!�AbK�O�o'��CD�qD�	D��<!~�U�$�|"�"�l"�,"�<"�"�\���������]"�J"�{D��D�D���������	�ӻMI��D�mD��D�D�-D�MD�ͦ!����D�}$ƝD�=D�]D�o��;�����{����	�[LI��D���'��'��g������MC�c��*�6��g"�/D�D����׉�7��������S�)���!�	�o"�c��OÉ�+��s(��L`�$e���\şkC��ND��1�s�<!�v73?���;%�[�2�ucjsI���(��*�?��x���H�D�B"~7"~.?��ߝ�߃���/�W������D�r"~"� "� "�@��5�_Eį!1Z��v"���o&�W�mD|H�?�S�����G�G�>"���?�4�f<���1#L�G��~">Hć��">J�����LI��D�iD�"�D"�"�$"�d��|�0��%�/#1.$�/!�/"��#�/ �/&�/%����gԘ�����W�?$�%�D�_c�4�����_�?'�E�����������%;k�_{�)���������������4��c<�O�/���/�����$�_ �_"���k�7%�����#��J�����;��i������ϳ����!� �?!�?#�$�"�?��o7#��&���JQ�yE(�BLm��W��+1��&N��*"~�Q�	̛��̛���G�ϛ��ͫE����Ϋ��_jJ��"��&���=���D�2���x�$�H�:"����'�"�W�"���?8O��a�s��'�7�^"���_G�w�kMC|���E�H�"�����x�'�7���yB|�#�$�X"~;���$⇈��D�6�1������I�Ӊ�o�g���g�g��	��mJ�K����6�-"�
"�r"�;�!�㉿������	�3"��D��D�����������GMI��D�]D���!�� �K���4���x�"�$1~O�?N�?F�?L�?J������$O���ݔ���������������i��x��!�?"1�'��E��������!�n�_����_��ϟ���P��VLm��/�D�%��É�_�ϯ@1�a�](��r��|'�?��?E����Ο�/��MI�"~7"~?���O��%�癅��3�'~���؇�ߏ���'�7�/�?�W�?�ޔķ�D�*"~%���o&�1�����?��8���:����@�N�Aį��o5%�a"���?��?���A"�/s��K|���o#�w���� �'⇈��D�	D��D��Z���=�kC�R���j��?�jÛjc���M�lZ�:,f������o��� ��(��L�9"8݅�F'����i���6i�+P72DE�­8PAq�['��_Q���~�������=X}���{��}���^����J�m�����o���ʗ��L*a�C��խ��|���ӷ�o����%��b ��֍4r5�2r-6�2,v���N��,��ܾ����e��>�ĬST4Y�&�ժ1W̱Ս8������9��o))���o׷!�Qf�m�Qs׉%=�k5w��5w3j�V��MX�-R�a���p�sG�{p?i�|�k����^k��e�1�Ã�}��
A��K�"��QPk�
�T�M�
���j��f�U0[��Tl�|c��{kᤦ�l�6�4Yl��ꌕzq�+�6���[f�M_g�MVAo�4��i/����b��%T�̠��7��V����@9,�e��Q�Y��6��6��*����E�y���jR�	�,�-����>���C�������ޒ�J|�럠dW���:r'�4�)�]�ή�S�ہ~�?�K�T8�*m)N��
�U��dp���Ŋ7�j��5��H);�_�q�^���k�$A�+���m]�<�l�=��ֶ��$Ԙm�����:�6S�����9)� ,��^Ycl�
̭�h�b9���2�`�X������i��s��N�����E��W8����O�4��%�|��.�o��I;�b�-l�����:� �S���y�U�?W��#iY����������l_JEl�=���N��k��=^�)��jˎ�*U�X�SS}�A�/��`�Q�&��y.k��׸X̧n�|�S��-����*[~d���	���9ն�lG&��s:��z$�t����9�Q�5����Ͷcy���:�Ь@���d���d�o;5���l;�0M����x���e���~�G:�x�qM�`'߅�|��ޠ@�k��ۖ]��d+��K/h������,�vBh;�̳��I?ũk�V�<���ʨ��j�����Z�ǃ���`O��H�ˣ��q�i?�����Js�����F������E���b��6
�=W��j�o�T)P;5����x�U'��Jݫ#��)XG�nב�7��cRS�9U�׮!ۤV�kH+����r�s��tT�m]sr��`�h-E����mbmض������m�zSU�X}�o�26�+��&��� ���jˊ�2���"�[[��l�L�2��{�$F�w:���w�x=GF���*���&e�
]40َ����V�`�vvk0�6\�=�zŹ6���� ��>Wh/�,H���'�Ү�O�e��u�f�;6�-v�ob���"@�:�S�w����ڶ2�I��aI��R��j�����m�{�L��t����Z�G���M�:ڗje��T��N��]�=�i�fK�cm�.�@%?%�(��M�N<B�8���t�{�}�
~ѾY����:l�S�v!�{fy�a��N_����js+M\�`i���)�}���-����E}찼���8�3�I��Y%��*Ѷ��f�U�f�ci/O����ssbia�s��8$�o��G��}r�e����vs���a�;P,�o�� �S]&E~��Q����lt.M?:�"�I1��N��Ρ�FgQD��y�h9z��7�ng�g�ģ+F0��B=�Vj�L
�,
l��B���]������r)�
�ě!���o��Fn��e/�\�_�0.���!�B�_��C�E	ğ��&.�o�����/����_ɍ����o����M+����C�����7�E��\��C�6�����!�n���^�.�	a<�/@�n�⟃�=�"�?��p)����߅�w ~?Ŀ��s#~{�_B�A�����B�W ⿃� �k���rp��Gi���I�������� �on���\�� �x� 
cL_*`L �2��Ԙ^��>ؘ� Z�1��"~8�����ɘ�(�1�RicΠ�ƜN���"~���ŏ���#� >�C >�#!>�C�"��g�.>��!>	�'C|*�'C|
7�'����#�!^�9��_�*?�/.��B�� ��k � ��܈/g/��"�&�_ �� ���χ�f���E�7\�_	� ~)�_
�+ ~�/�F����_	��U�_��!~#�o��k!~�Jď
�R�=/��	�w@������F����?�O!��!~�?�B�v��wB�cj?�K�{!���_���!�U���/��>��0>��O!�c���B�'����#_�R�!�?�?A���+���p#�{�����CzP!�T@H7
%�����C|(�
!�;�U��Q��(>d(M2�"	H1�Si!C(��AQ�`^ć2���Q�L�?�Ϣ�
9�G@��?�V6d�Z�_ȥ�x�O����q���^|
�g"�)?�B|*ħC|�O���N�'V���B�;`_���H�R)�YBfRa!�X�N�'M���}!���/��i͙Ps��z,�������:q�
]��P-M���b��b��Ť��:5��8��?��YJ3�,Sh@����bP\�;���!ތho(�qˤ���y�F�iyCىs��uI5��6C������(5#U���v�6��[�<���È!ҀL'ƈs!w ��8�Kܓ��d{�A=�xhT�`!�8�S�G�POb1�����b�dR�y�d��3矼�&����fk�;�}4K��TXțX�[��V\����>�q�<mȗ4S�W
=O�	j� j�c�ħ��V�c�CM�.��,m�W�q�V��@G��� ��,J<@��eR�7�p�����>4�"	I1��C�����BGQD��yi
=���Q#P�8�8t"�B)��xZ��
?t<�@!�N���UI�g�S\�ρ�\���� >�3!>��S؋/�x=�:�/��_
�!��g�E�=\��@��M_�o��n��a/~�_�0·�� ��?�σ�!�b�_�AC��!n9R�~�o7�.�n�~��߲.�B��,��Sa���ص�4��~��h���z���P�e'o�	�[vBxˎA�P��4�̖*�E���F{�e��]4�dY��4S�N���C��A�Q���nӽ�wф:�����~�m���f+j�MC��n	�6UfA_�K[�+�/�C��(��Y��@�ot�E?T|�y�[�o||�n*i�����i?8�fP7U��h�ѥtn�U5�D5��e�P�溍��p]yb�����A�}C%����2�wD�����]�|3��m����g��9m{<K���k�L��Lc�d]-#YE�%�y���T�+��H�Jv��4ׇ��h�6LwI�g�g���Ao�̫�d��J��չEvK1
��u��l�8g�J%�j9�p:r��]3���!3l�B[���Z�q:����b��W�ޖ�N��IFҮ����uN�绷�0E�9]0%7O��J.��LOD��57r�M����t�μ.JF�d�ۣPΔ=yhlқf�#7�H�~u&���*���	�w�	n'���vۥ�AGY����^A�5w�V�Q�Y�f����}��$�.?-=-?-;%MW0#W����î������b7�}���)��G�&������� %��㺒n���^�I�sC��;Z1���q�<�a���tc���ΌT�	j�nm���O���M��m��l�Ҷ?9*��h��E�/��m����_S]����_���!uz�f���D��U����-�Ϋ��Y�E:��`i2�|H?[&p��l�r���>[
�>��M��G˿Ns-�X�	�,�\,>z�(j1V��8�r�D�IBlue����ds���[e�F�{&��֯��ۿ.J���^һ�t�I��3����E��s�E��Bg��5ӳ�)}�#�S�ӧ������R��m���u~��C����ۅCo��a�rsor�����@U�'9�Nr(�ɑ!�]�)�?O���}^�g'-�vNZ�;}��r7-�ӥsfv������ovޒ�r2�r��錆M�,�;����*��N������e�[�Jy?m+e���6�*!�7��d,�:���&k����>gl�<����ݜU����b���Q#�f��I�]��kE6Pۇ�Qɬ�����l����<�.#s�dh��)s����U2_��o�1���OIs}<��7/z���ؤl���"NsN���)���T��R̙.�^���]&�Z�Z��Wd������R��l���6�Q�����B�ҥ�Z`����Te�b�y^$c�Q���#uIȰ�R�5FA_�&w�@�P���0@d�q��*n��cL���H��&���4�`���ߺ�Mp�l�uo�ܛ�c�9nYn�Rns�(PW�͉�7'��Ȑ*���bl��I��3EzFv�Ɓ��x�m���'a�75�r[���H�PPk�:?"�[�Ɏk'��w/frkͬ��ֻ�{�8�]28�Tx �O�e=�ًf��C�E�b#�W�vn<A��Z��߶����4�4�`$f�<EL�cFA���Z�Z*ө��i�fK�cm�.�?6���\�Q#O�B�; 8���O�A��>8qp�˕�?U�G��4����I��b�,��"�(��
�(���Ѩ"���Fi��#�#�D�DZi�"�~d#)P��he#T2�Z�f.�/���	�_�K!~	�_ʍ�؋��7!���o��u%�o���!�
��kd���
�wA�m+��	�C�܈����� �I��(�?�A�6��C���Zħs)�U��_�� ��	�_�F���ſ� ���� ��B���!���D|D
����_ ��������#7�a/�O�8�a�CD�B�Q�?�S`Q>B��A�/���ϣ��A4}�`�$*�b�
�ҢR\Q(��`^�G�e.>�T�?a��gR(Q�i��N��4?�Ϣ��:]-�K���!>� >��B�8nć�?�3F*�O��4�O���O������.�τ�R�/��B����_�|��+!�a�@�����*���x#�υx�J�Gr)~1ğ��� �υ�����M��_
�k�
���WB�R�_� ~5�/S��Ӹ=�� ��B�5��7C�u܈����; ��q7����@������C�V���ǥ�g �Y��	�; ~�?�Os#�q��_������&���W �5���A��*q�K�_A����
�_B���7�?b/�G��?��+��� �'���C����Jć��Q|t/�>�7Eݝb��F�EP\�=(�螼���e.>:�&���1�
�>�B�J+=�L�E��O�����p)ﮍƻk����h��6ﮍƻk��ywm4�w�F��x��6ﮍƻk����h��6z<�'@<�]��w׆��R<�]�w�F�ݵ�xwm4�]�w�Fs���h�ﮍ.�x��6ﮍƻk����h��6������r�W˻k���R���w�F�ݵ�xwm4�]�ͻk�ٿ�6z��ݵ�xwm4�]}��ݵ�xwm4�]�w�F��ݵ�I|�b.ů��9į��+!~�_����؋��oC7B�-�o�� �f���W���)\����� �A��A��܈�����!�E������!~�?�!��F%���p)~?� ��@���>Ŀ��q#�M�⿀����⿁�/!�k��⿇��T">��������'���C�����1?�'M<6��ۇ
۟BۗVjl �?�76��06�Vvl/����£��g��c�S$cO�ǞB���P\cO��ƞ΋��'�?�F�GB|8ď��P����(�Q���\�O��4��� >� >����gA|�ȃ��χ�l�υx-�B|�Jć�ȥ�����J����j���x7�u��7@|3� ~>�7A|#�[!~�/�x�J�G��R�
�_	�B��_�K!~7�/b/�
��al��M�_	� �j���׫E|����{ ������;!~+7�oa/�a�߉0�C���8�?�A���U���׸�:����!�%��_��W������ �3��!��A�����B�~���ƥ�_!����!���	��F�w���E��Na����S(�|!�o�?J����u��T">b�������H�S��Pi�S\�RD��"~\��ǝ�#��?�Ϥ�������� �Z�qg�D|X4��� >��A�X��1ˍ�H��!~:�H�����)��S!~ħ�D|D��gA|ė@|1ėB���ɍ���oBF����9_�?��!�F-�r)�|�� �A�B�?�υ��܈��^�2��a���5�/������B�
��o�j#����A�f���@��܈��^�V�a��@�}����C���Jć��R�s�<�?�OA�����F���ſ
�� �7 �-��_�����߆��U">|&��@�7���_C���7��ob&�g��a������ ��?�C���J�G<����>4}L_�$�'�ӃJ��Mq�PD1�x��\|� �8�T�1�
�A(1'�J���c�R`1'S1����Q����\���p�� >��@|���}����ً����#�'B|"ď��x�� � >��x���h�D�&��Kc5T��_")�4�f���3df����9Jۭ�v*!�Yizz��1Y�Ҵ1S�;��^Y�0&��[֋�b�h��*,&�͖¾�I���v�C��w�CV:|����*1Rz�ˏ /��:���-ˢ�vY�Z��F�u�QF��Kz���f��uS���B��X�\CÜ��>wt���@�=�Æ�o�cj���0�n%�͑Z�e��� Mv�wF�(X�-��wF%���ȘE4S̹b�����)�y�p84��|��
�M5�Җ�T����[Ŷ� �SuI���ط�6o	[փ�Y��Z�w� X�M�SͶ.р�m��ws���n&}�A�۠vܺ��Y)g�a6Fl���fw^d�9�k�G|=� }ЮK�}�fO7�۰Q܁��V,�v1�6���	|�4�]e��"�f�z�m��ߎ�\̠o��ن�z�*J>�덷�t⍷���bV���n�~R�h[ξ;����V��9|խ�ȿ��Დ]�?Mۍ"�9�u��J����b}(�X_n����3����K��0b���؁J� Z��~~l L!�����߉��Fq���K���y��>v��G��3h��TX����Kzi�5��F�1���&��d�Z5�9��iT�l�w/�c�<��X�\j.����@����~q)AS���f�`�/�,����Dت�k��?j���Ro��++EI���&#Kc�"*17,�Y���\%]`u�!�_Y�y4Sl�Bm��V a�!,��6�Um��2m���6m=��l�I�L�<C��-�MSm[
j�����X�m��-�N,�v��M�ms������͚*C��d4�ض�`��i��뚤��mzǥ�h����f��XQg�f������T�U��*cu�����!&���X�yҡ�C<Ӓ�⡎���y���m�pT��ZC�Z��Rd��q��r�r{ʨ�EΕ�������݀c�a�٤D��#���J�l�{���jU�8׶3�o�T��q`;9v/O~2�t�s�F#O�L��_�� ���ί5��Y�EPcmjh0[l�YcM�*�C�Ղ�N�ln� @�\&�A���W��2�5FSv��[���~���"4��8��Zz�P%���d��J�1.}zg��q�/M��͹��Zce��l�k������C��� �o�����-~�J�ݚ�ZC�ܖ�l9W���j9�vZ��F�V��ՙ��Hi�����tX5�z���}f�2����۾�0�i���)q�Yw,c��z>�ZDgN�˨�����'�R�)|�n���wu�f���
������{N2o0�s|�x�.o*�����(tS)�O�e�j��đ��J��T�&�v�o*�>F��:��$9̢ĝ�~.�"�NR��<�I?��?�"�B1�O��ƧS\�S)��i��I?���ѝ��4����
_L��/���G��R`�(��%����U�!:�.�ρ��_��7B|��r#���x+ğ�0�C�B�_ ��σ�f�_�Mj_���� ~5�/��e�
�W@�Jn�/a/~�oA� ~3�_�!�j��⯃���"�=.����C�]�����!�n���^�c�a<	�OA����O@�N��W���\���A�k�*Ŀ�C�^nĿ�^��%���?��O!�C���?��/ �#��_ĥ�� �w�������+��F�A����qF�?׃B��F+�C���Q`q�)�����q�j� ���N���N�H�S�q����aW��(n(/��07�� ��!~ğ�# �,�	�!��z��>B�שH�{��x�o\�w��ƅ�˺�C�č����a������].�Ve޸4����K��n��n�P7Ӱ��N��|�'����'�ݽ9-���Ԯ{�(�4S\�B=n��!�"t����m����A�[��V٧v�f=�qkm6Uꬂ^h�����ûRg�z0ĉ�=�>p�?���Wzԥ��Y�	ͦ��ʨ�5Ε5ȳ��t���'[�V�<�@�yƪed�MJy+��aQl�5GF�T���|E�ɗQF��Sg��w���<�!#c522��:�� ���*�׈��y���Xj�-��o�%g�qa��t���	?�E| ��P����4K|0�k|/���>]]��z�:H[�
:v�hq��C���Ƕ��4}�L�$��b�/���K(��"�(������<�oFm��4q�\�QM�)��Z��J
?�@���R�she�Tr7'��~���B�b�_ ��!~�7C�Bn���/���c9į��)�/����/U��w��⯇�k ~�_��B�fn�od/�v��a���B���o��{ �>��S-��q)~�?�; �I��wB�S܈��^�K�a��o@���2Ŀ
�{!�M�E-��R����
�@���΍�ً?�#�_ �0��
�?B�������"��^Y	4}B/�$�Ř�O�%����SD	=x���\|� �8�d�1�
HF�$��J��Q`	C)���he�E�.ŏ���?�φ��?�Gq#~{�c!~��	�� >��!>�c:������;1!Ż���#�HB͒0�
K���NS�w"ϣ�&��n�ń"OkN��ӣ�fc���8(9I�GM��1T�5,b��]�۾���h��M��Z����Ę��fJhV�c�4��4�v;1��o:��}1A�����0��/�ŕ9�e�jP�m�-��e6�05O'w̱6��IN������D~3a�^�Q_� ���t���.=~�8Wן^�.���n嫗�/��_��Ί�	.u�S��	�V�>��۱e�[��YvSa	�b��w�&��.�m�)����$�EM���x5�F���>��t���%�Ǻ��5���Ow�I��*��~GM��
%�J�'�F�$�D1&��O��O����K�P�`�oF�B�g�ĉ�c4�J�$���J<��OE�%�P�a���#U��p?��'C|�'B|�O��	?���ًπ�|������ >�s >⧫E�.�WB|�� ~6�W@|9��_�^|�7!���B|#��C��-/@�I=#$.�n�|�oYJ��,�Qa��c��F H\��V��U���z��F�͕X�N���>z�,~�~��%u��>��)�^�Z�� ����vp����$�ߋ�Qv��F�l�v��
Aq�A���J��A�m+ǰ�8��)7�Ů�'����}�����-��l�2X�T�����u�0ϟzN|�u�����V���X=��(#Y�:%���J�Ս���2n%��L��}���
����Z�\C�8Ѕ�M��O܄��L\�}�A'�N�XHF�d�v1A�Μ������Ygd4�
���s��(��x�4��7Bɜ��Ns�n�2��5�z5��wd1����n@+V%���zq�Vmd�C3�P6�9e�١1���1ڄsչi�6Zu�����MW93!g.ߏ9��\=�6���.P��d�^�3�&n�{��[V̄�h�	Sa��N��5|��f�	��Lv+��g�Ө�P+O�Vvu��5|��u���s�ˤȿ1<!����h��(��})Ɖ}������~�������p�э�'���#�S���
e�i�RO��'�B�M<�B�x������+Ąb.�GC�X���0�������F���!>aL���O��	?	�!>�'�D|�_\�/��b�χ�<�/�x-�p#>��x��"�J����*�/��
�7@|��U"~¹\�o������/��y?����_�+ƥ��B����A�
��D%���R���⯂���_�%{�@�=������[!�v��
�wC�m*?Aå����?��!~�?�Or#����@�^��2Ŀ�@��Ŀ
�C��j�ƥ�� �s���?��O!�c�������B?B�/���!�g���P��ĝ<��ԝ��ԃ"��u��C�M�FqM�&�s#�o��'���'�0&S�S(��JM
��'��&�&�������R�H��gB��?�ς��y?I�^|$��#�q?�c >
��B|,��A|�Zį�R�t�τ�)��� ~*�gp#>����/C%_
�3 ��!~&�ς�"���åxě!~�!���B|7�ً�� �Eğ� ~!�/���!�Y-��s)�r�_�A�*�_�!~7◳�	�oB�A��⯁��=���תD|�\��A�}/�?��C�܈����'!�y��4�?� ~�?��@�s����jy�'��a����a��߲��Nz�f���
���}S�axjy�g��a�Ǟ���ܷ�����o:9H���Ǡ3��L��S#,K}�Fkh'Ŷ��~4�d�Fk��W�N�x��<�a��Z��hb/eGk���m3ZCo���75T�a��#,�n>�2y`����j������H�h�0�t�ʹFS���T_�j����Q���%������t+w��֙�8Bǩ�?�����::>�&}�]��pPp,Q�����C.2��m���iH�l�i�� �OKO�O�NI��ȕ�����z���P�&��6����K�H���~k\�dб�p��n���^�I�sC��;Z���_�Uy�ÂO/l�R�8$�u�8�MJ?��O6�_,@Ӻ�O"��2�4��忦�:�ӿ�H�?"B���:y���3Vy4�<}]�A���!◐Ȑ�*�p����c�y��:��H�?,M���g������_����gK��G�����O��h��i�E�5��E���˭EQ�CB#��8�r�D�IB�'�_���<���G��C#�5E˿�_�pQ>dR��s��$U��5y��nț'��*�~.P'�2�M�0.��/&_�6�Q�|�f�zW�����b��e�2<e�Fʶ*��a��˛��Cr�5����y�))6Qv�]v�]rvi�|�m��u�UM��Ս�i�y�1J�gv�	i�V����τ�;h���`8'�h���SՉ��+���f����X�%c�ȤA�Y�|�Me[p�ڳ6_o1�m`ϥ0�������B�K){���>䷨'%�,I���xZlRb��;.ۈ��h��l�F�I��Z�E�LA�dt��sB��c���Q�t��0�C�p��]���x�����O�H�$��:]N�%����������kP�j�oF]�����I�#�����[)���i�����n���n��n��M�A%��&_ť�� ~;�o��� �Q���F�������������g �9���/B��*�t6��?��!�]��;��߃�������/!� ��⿇�o!�+�? ��A���J�O^¥��4}����?!������F����'���(��T@r ��܏V*���܇K�O!$��&�V���<�O�#(���(��S���3(���)�d/�Of/~ďE���a	����I�������!>�!>��؋φ�b�������σ��/��\���<�K�o��*�����7@|57��ًo����	�@�<��@� ��!��j¥���
�B����A�rn�_�^���a\��@����7B�&���7x[����'r)������; �n��
�w��^��8$Η|뱷��}��~�x��.��$����}�������>vb�x���{�7���WO���{�����u{<�U�%�u*,�,�������y�����������Ps�c�_v���c=�u��}L�]Zii�����i��z�7��h�t�J�2�h��^��d���C������P�xj.�^���uٺ�c�z��[d�K��A�y�8���\�)L?�ĉח�?Λ���R���q^��Ö�Bϔ��*qI'��,q�S����3�;+�͋)��ɋ�8yn��u3y��LF'��u���ʥL\��rr��MG����
j��#4m�ő��gh�=��{��H�����qs'���F&�j���R�8����Z�K�֊�A�� ͒��
Ky �}��O6�>��f��i��gi���z�!e'jb7jbj��?� �D�CM8l']O2t�G�m��}�A��x�QI�A�|ޡ����G1e��WR�����Ijo�1���ڏ�J�C����bj�oFwLR��ĩ��RO�PRO��JF᧞L���J!��N+�z�Jdp)>� >�C >�� >��؋����1� ~�'@��������\�/��B�υ���B|��s#>���2��Fz����
����_	��שE�Y\��� �
�����7q#��^��a\�K!~	�_�C����/R���\����@��_�WC�F�����؋�	��B�A��;���B���oQ����s)�I���A����o����|���nc/�y�a��@�K��_���!�U��Ӊ�~��z�����w{���i�-��8��%�#*,u?�a'{�I߹����w{��~�i����;������ӽ�:���`�&�z�G;K�dG���4SZ?�:����Y�i]�z���v;��~�G�����~�Pʾ�cj�M��X���-��N�57YX�+����[�ib�"C1���*��ёu�[�:k������~?����e��s�4ϺG� �ee�WU�7���L�__�
��C�ȡ�#� ��5Q�\)���̉K�M�\	>C��]��"������zs�I`��%�'0m�B���sshm��a���2�Q�[X/Es֟M�6R�\���9�v���Ұ���2r�Q*W���͕��'C0�[ufA��Y��(i�;����%���w����٤�J��պ-����U2rU�+ϟ�P2W�S���u�����O)aJ�����a��fʕ�)$e�"(���lre���Ŋ�j��[c���A��M��b&�KP$c�8�[�&[WP���ۯuΖ:�[�O�)��A�"^4�{۱�i�����+��Q�w�7���<�7H)$eva�)I�����`tZA/4Y���B�r�jl�\5�0�M1c�(i����B�u��x��J�"YS�P)�t7��r���b�^d���,Ӛd������n�G�^Dj[��xl��;�>�K����������}T��,��u�H!)sT{[�\	>����I�j�V������Ɓm�"����t�lm=+`�8���Tg�l���d�rʖ�=xx����8C���8]<�Vs��-u?wS�՘;�R7���:�6�5W��ɕ�r�z&���13�Ies��M�V�p��)W�T�J��j��7�	��&��`�l��ʪ��Y�~���u���M�6S�\w�BRd��4*I���a�_�[�hK�Pl�74��DNOd��j�K�s}��Jj�;�{a�2�&qsd$N�%�'��U_g��v!���)�3m���?�d˃V��l��l�q��S��5r��h�"���4�}ORH�*#NRr#���,�Pkfԋ��eMis���CfO�7�7�H�󦨞^qlru���2B��r���Ja��BR�+�g�V0[����(0} ���MU�N�h[O\��2�7Y��7�B6ٺF�vZ��v�����A�����V69�1���*u�l�T�����ƹ@��9O���팕����0�\��l��0.r��2�iMJbi*k���._/0�������Ի�H�|���_nj�����ZJ����;�BwF���B6���r��I�*���V���bʕ;3eZ��%mR6W[��j��\)�x-.�n�re;�hy�T�r��)m����I���Ff����*7�\��S�`ϥ�H���?�M�h�%#�
�E��#۹�R>��rm|��o;��	񆊌D�)c��.�P��Z��Z�A������*��k�ui]o�h�zK�o�0h0����w������� �Ki��eI��c�ETZƥW�%Q�)�i�q��7�>3���W#�+����J�zZ���)��+(��B�U��뤴�!m�7s)�N��
�B�-���s#�F����'�#����� �a����m*��؁j�
Ŀ
�/@���_�����{�oC���}����C�;�� �A��j�Υ�� �g��⿃�!��?ȍ����AO�CS�| ���������4_�?��)<��6���6�"�H1N�O�M���QD��"~Z�⧝�g!ď�P��A+5�T
��ش�&���T">�?��c >� >��A|4ď�F|{� ~*�H��t�O�����i?��"^å�?�!� �K �⋹��^|��E�o�����x��B���R���B.ş�!~�χ�E���/���W#���
�W@����WB�e�T%��J��⯇�k ~�_��B�fn�od/�v��a���B���o��{ �>��S%�����]����'!�i��	�Oq#~;{�/A�>��Ŀ�C���*���7!����8̥�/!�+���?��/ �3������G�@�a������!����?�D|�8�O����H�w���Si�{R\ӻSD�{�"~�s�����OF�����(��Ch��S��Q`ӇR�O���>P%�,�R����s �l��#!~7�G�?�' ��� �q?�c!>�!>F%��r)>�s ~�g@|�O��Lnħ�_����gC�,�/���_�:����S�p)��-_�u� �&�7s#��^�B��a��B����C�ğ��p)�J�_�k!~�_�C�:nįb/~3�ߊ0n���!�F��⯇�� ��ߢ��\����!�����m܈����� ���,���� �i�⟇�=�K%�Vq)�}���oC�[�Ŀ��r#���?������-���/ �+��⿃�/U">���ɿ!���������?!�7�3�ك&��02{S��(��>�R�=)��^Xf_
!�?�lf�Jćm�Q|����<�"�<�b�Di��S\��RD���">s{� >
a�B|ćA�h���p����1*�n�R|
ħB�$����?⓸��^|&�"�\��B|�gA|��C|�g�D|��\�������x=� �⫸?��x3�/@V����7@�� ~>�7�D|�b.�/����/��e)�/�F���ů��k����7B��⯂�M�J�O�̥�� �n���o�����ɍ��ً��;�c��o���!�Q�⟄�GT">� ��_���!�%��_���!�n��f/�]��a| �C������� ��_%��n�R�/�+��� �g����F��������!��T@�����A�?X�/�����D|D�g�鳆P$Y(Ƭ *-kŕLe�E|V?��N��s�p�?�G�Je�N�g��gB�ٴ�Y���:�K��!>��B|4��B�8���F|{�I?a�A�T�O��d�O��)��)*6�K�?�!��gB|	���F����*��G�?�o�����u_��G�ğ�!��C�"�?���؋_
�k�J�_� ~į��� ~�/W��.��g� �7B�f��⯇�� ~7�f/�N�a���C������� ���K%⧬�R����?�;!���wq#�	��_����^���o@���:Ŀ	�oA�k*����!� ��A�W��ɍ��ً�	��@� �w�?�?C���������i\��d����P$�=(���TZv/�+�'E����l?����٧ ��T@��J�0Z��A~�
,�$
!+�=X%�3�q)>�� ~ď����c�{�1?	a�C��O��X����D����U"~J�o�R��\�σ�L���9���܈��^���@e_�!~&�ςx��!�T%��s�o�x��o�x�7@|#7��.�/A@��!�/���!�"����S���.�o�����/����_ɍ����o����M+����C�����7�E<�c�e?��!~�?�B���7��g/~Ŀ�0��� ~7�?��A���U�����X��?��!�]���C�{�>7����%�D�@���-�� �;���V���\�?J���@�������� �on���\|N M�3����K�R(9�h�rzQ�9}(���BN�lNo��O�Q|�p�A��F1�J��Aq�N�hx�s2{�c ~,���(�������H����P���̥�4�O��$�����)܈��^|6�#�|�/�x-��@|�@|��D���\���x#�WA|%��@�⫹_�^|#�/DM� ��A������oU������WA�R���W@�2�_΍��ً��7#�� �����C�F����B����R̥�{ �^������!~+��ō�[ً�B�C�������$����T">|���B��
Ŀ�C���7�_`/�}��a|�B����?��O �3��@-�|�_�!�?�?A���+���p#�{�����s{P��T@n7
%�����s}(�\
!�;�U�������s�Q$�)��`*-wŕ;�"�̋��@��s5?
a�	��@�Y�R�g@��?�G���W����\��������q�?��Q�ŧ@|&�� ~*ħB|:�g@�t�OS���}\�/���?�K ~�τ�Rn��_�f�1��!~.��@��� ��j*��/��!�\�_��C�b�?��؋_���e��WC�
�_�k �r�_��Swr)�&���@�u#�_�7p#�����m�>�����!�^� ���{T">��g�r�����⟆�� ����;؋��EoB����_��7 �-����D|�.���B������� �k���_���A�A��;��
�!�� �O�?�V��{H��Q"���M��R0�Ms�F�5h����a�L��������V�o;���4}�s,V�4m��T�b��+�[;e�;'ܧo��b��ܣ��b�R��֍�@������z�b�zIa_�$z�R;�!��;�!+�_��]<)>i��G���b��O��eE��#����b�6ʬ��2�f�X�г�U7y�<��SQ7��nN�b�wpsf?4\����>ڏ6�RM��p�nߖŘ�B��,(��g��G	Zǘi�����C+�`M��$����f�#6-%�ℜ捣��QY�t��B ��p@����p�H���p1�%z�����J�Tc�F�Zbl]���4�ͺD�1K�uIԥT���\fK6m;g��� �hP;F�������E$���#nlA�;�t��{K}�m�A�񡭠%��b�R���/�V8�%��#�!
Z���[疪um����p׺�pK���E)�G,�tC���B����iC�����P৲wN�:�n�s
l���8���t��ͨc�pxȞ,O�d�Ă:1�N�J���T'��e�Zv9Ԅ�+��T��]K�q�ÉGH����N(�ط���[v�����~e
6g1��{fy�a��N[}�����+,>��]�h���	�W:�2�P��˻�_��?s�����aG�����@{��EƖ����gƾ�q���ߏڿ���4�@?�_����^~�X��<�O�����y�<^��=L��=B��=�u��J��Fq�=H�=�K�T�=�ߌ.��v��y{�3T@��J޳�RyOQ�y�(���(��ݴ�yOwpyn��{�o�v����W�{�����7i������7��}����/�c�C�J/�?��e�Ǟ���ͷ�����o:y.�IN��
�K���h2T�Ԛ���U�ۗ=����=�EHg/̓���ti��K3��)ui�͒�8� ��Ǻ4�\k��<OK��Ks�S��K� �C]�.i�ͥy�����-ͪ�2������U�xa��Uz��`�J[ �_����<����ܭ��#�VN�v5U#��Fz���b4n�j��*��`�&�ՙ���$l��2a��	�9�	�+&,I,�p�h���t�U�q͕��L��HIӲIU��T�vJ��eǟU��RώU��\58���>Kٳ����?�ɿ�fɿ�
˿�]�Nӫ���;}N����4S��\�ע&�BM�AM\�H�k���h]�����8��\�tT]��(����eR�7��g�������1zb��X'����������܌���~��|������1zb>FO����=1�'�c��|�������gs)�'j} ��	�'�c��|��������GO�b�D-FO�b�D-FO�b�D-FO�b�D-FO�b�D�ZFO�ɣx-FO�b�D-FO�b�D-FO�b�D-7�'jُ����Z�����Z�����Z�����Z�����x������]����Z����������=Q���Z��'j1z��'j1z��'j����=Q���=Q�������=Q���=Q���=Q���Z��'j1z��'j1z�v�c�D-FO�b�D-FO�b�D�ZFȌ�R<FO�b�D-FO�b�D-FO�b�D-7�'jُ����Z����
⯁x�����Z�����Z�������]���*H]���x����F�v�n��������f��I�io�b�P�����Y�]���x����!O��I��N��X�Nw�l�I1��,��A�&��������N��'$�h�y�_�D�-�}�fҾ�Po!���>|셏7��-dKq�^�W��]�v�iŎ���:���3$����+���m]b'���6�*uVA/4�����=2��j��U�;��Xl<�#�����/X�ۣ�Cz�u��"�/���%��B��suEy�����!C��A��&e2z�b'���X��Ph�c�/��
�q�W�g���dƂh7jOtFF������ũRZ��`Q哥m:�y�/9�>u���S��r����
+��b���_$��O˵���ö[v<�9!�Xh��B}�
�Q+M��:Ԋ��}��ib'?��p�n�C��Z�"iTA�#���T)���;����G����Q���
�����H
�:=B�<Nq<Fl�	����Ī	��9���U��P�2�R�"�T��~�
��%
��Zق�*�iQ�~-�]���	���:��A��!7��a/� ���0���!���⿃��������(�Џ�/���NSi���"*��F�������Q��T@a0�RD+Uؗ�/�O��
���S�x�.ş�gS$�gP���?��*�#x_x*{�a�0� ~�GC|8�GB�X������/ĥ������S >�ӹo�L|��D�_�E��_�3 ^��q\���u_��?�k!�ȍ�J���_�0@�"�o��&���!�\���A�#W��PWy�KR����Tx����V���4K�J*�p�B�.I��F�1���&��d�Z5�9���Ve��«��a�p��5�5wj�:,��NwX
��6JM6]�����#�R�4S�c
�O*|���!٣���a�$�/eF3�C]����S��7r�2�D
��#�t���
���=��S�D�xu^T���kI,�m��䗒�&Csed�'�����'�JQ��)*�SS��-����*�<��VԦ�g=���S�$A�W��w2M�c�< �Q�w���M��ON���\r8Ar�f���s�x6&~�5���Op���W20y�w�mp��r�9۹b|��&�e�\��0�KF7��4�$7M�J��O��Zi1��>�d賢9N��=�-Q
_$�m�-모�<���*�h1-����wMl<�>+ZC3�U�;b�
��:��r����wGl���k��r��@�I�g�7<��)z��/z�")z�b,�K��Eq�I���Nѫ�ߌ��}L@�SE_Q(E_�J}B�}F�}I!}M+[��J�Z�p)����c�A��A�o�;7�f.�؏&.�Ca���{Q(�=i���)���Xq �PܛV���J�~ģ��Sh��S)��ac�P*�q�D�̋��A�ş�acć@�h�?�GB����sT"�h��'A�d�O��x���?����O��<��	�9��?�!>⧩E<���+ ��gC|��!^��܈��^�\���-� �uo��F��B|�Zğͥ�%)�_�@�%�_̍x���į���cį��+ ~�_�WB��_��?q)�v���o��� �6���o�F��������6���� �!����U"�ȏK�/A���⟇�!~Ŀ���g؋��"�w!~?Ŀ�oA�;�>� �ow�ü���şy�/y��o[-��V���⯱�o�Kި��-��no��C���ߨܚ.�������m=������ �Vr4K�G��}�D�'^2�f*�P?� ��d�kI A(p�~�1�G{�ĥz�x�(��x�R��l]R5�M?������cN/s���g7���L%ⁿ�=���@bı�U�q�$z�{�q��*z+IdYYb�c�=����tߑK���Sa%9Xl^;��|�Ǵc�6zү*���c�Ϲ�WU��Q�P���Y��*�I)�L�~U1�j�a��o���.fT��b>�:��U9̢D�*�I��rQ��c�E	��J�VW����Օ���mu%ܴՕ�o�+A[]	��J�VW����Օ���mu%h�+A[]�Z��J��R<��J�VW����Օ���mu%ܴՕ�o�+A[]	��J�VW����Օ���mu%h�+A[]����X�k��V�}����J��VW�i[]	��J�VW������bœ]u�Օx����Ӷ��Օ�r�mu%�m�������5����-v3��L3�*�b7c �2�$Z�A�aF��f����N<Vfd����6-v=�pj�8����2�ꤐ:=̿:�f��n�'t��ސ1���7Č�ukW۷�XoH7���Z��w|(0��I�]�jF�s�|�c�l�����z��q|�=�/�T��b;�K�X̖,kM'��2���)O���<��
�ʹ}%��d��2�F�L\v\3�G<Vi�WR�:Tᮛ���m|�^���^ی=4ˌ������F.h�����x_�;l3��&>@M���x�k��Y�F.�:��w���L���3��~�LM?��d�)�L�6�t�k����x��0s��7��3G��3�F(03�B�F+5s4�?3��N!̌���9F%w�NI�R|
ħB�$����?⓸��^|&�"�\��B|�gA|��C|�g�D<���̬�����x=� �⫸?��x3�/@V����7@�� ~>�7�D�����]�r�_�K ��_�B�Rn�_�^�:��al���!~#�_��!�*���W�E��\������!�6��
�w@��܈����m�a<�O@�v�����!�I�D%��w+��_���!�%��_���!�n��f/�]��a| �C������� ��_%�gdq)����B��3���?q#�[���ĥ��Q*�ԏB)���� �
�ԗB(������wi/��-�a�-�Gi �R:�
+�����.=ͻ}CK��iݜ��9u3�=K�縥�ͮ縕�Z�H3�NP�Whi, L�@/�9n��;�*-A��q#�m�P7�l����Rq����ـ�k�CT�=b���B6�*,���dWu<u<_�.����f�I����P��,]%{P��.��"�2�t:���O���;(��ǰN�Ri�OP\��)���y�/�f���2��y���5��"P�
�R��T�n
��
��e
��UZ��=�yD�t��/��zz}�f)E���������G4K���e�W��͏���Q7�؟:��f?��l�2XtF�P/M��s���"|��<c�t�xB]���E3���u��n4ˬ�����IƬ��^��R���z�t����y����Υ'�]�>���b�h�j�u��Q�m��;�y��e<�9��Fǫt���gW�a��J��g��q�G��75T��+����r��N���SWb���H��#}��\�w��?��~���c��I��1�`_����s��^I�5.W2�y%}�[I7j�t�פ�YL�LO��Ѻ���/�J6H�D*�W�.m���̭=��$��Io���f��}q�����K������%ֻ�b�j�tFY,z��y�oU��vNY��)S�X��cM��&[u2�ݥJ`AS�2uʼ�[F�d<l=�yx��Ĺ��sw7�J�`�1[�-W�'�(#S{�2Չs�ӮU2g�ֹMl�%c�Y�;o��8�|�6X���a�N�/`�5����e�;g��X�aJ�_Kތ�Jv���~��Ԛ�>U���=O���#���6���z����N��K��iFY�B��>�P���5��%˒i��T*�,�[����$��i���`��,H�H�$�
h��B��I��V�Q+٨�������񧥛-��������J؎Yz��?�%l�c�R��ʶ[ʿꦫ��,Jt�8�eR�w�(��D�u4}���l��j*�l3�UvETv-/'�6�3�8QvM\v��J��C���E+Uv;�_v'Vv7�Pv/�l�*ybg��\��wA����?�; ~'7�c/�E�a�
�{!�5�	�_���!��Y-�?�R��%��C���)�ƍ�؋��C?C�!���B�O�+����"~'��g���gP$��)��~T����n���܈?�\�� �x�I��AT������R�P��R`��P�����V����q)~4ď���!�,���@�H^���^|4�'"�X�����?�c >� ~�Z�p)>�!>�B|&�O���܈Oc/��uc&ėA|)�C����!�D%�g�R|�7B|�υx3��C�����7C�Ec1�_ ��A�B�?�χ�!~�Z��ť�+ �J�_�!~į��˹����k!��q=���7@�f���7B���Z�_ʥ��!�� ���m� �?č�{؋�	�{�3�<�?�OA�.��wC��jť�� �}���A���6ĿÍ������!�� ����?��/!� ��_�E�^.���C��A������?���x]w�Xן����t})]oZ)]
_@���P�~����*��e{��t�^��Ht�Qw2��;��ҝB�N�E�n({�#!>a�@|8ćB�(��a�U"~��\�O����� >	�'A�dn�ǳ?�F��C|.�gB|6��A��:�D�&��X[��i���֠�6[�&6i��2���)����0%�b�oY}Xu�4���
��X�RÔ�U�0%:�w�)��yZ7M����y������R����KK�렡��H�*MvbN�[M3��(48�n9<\��aE����>f���7,�n����Dz�[����;�e�Q�m�#��Ԁ<��V��'׏����UV��tή�#����<�$ G�(#�M}��U��s}UyV_���*x�[����]R��������0��~�z�H�a�[ؤL�S���LY������:��t���[]6��0���Yy�A|Բ3�ӲQf�MB-��a`*������qd�P~�s�y�+%S�;�ha�I�x��<N��d��ֱvX���֯����j�Y��&�`����
�Q3�H[�:��3E<��0�V�1�N��y�nI�w���rP~1�R��
+��[~I;�t�-eRq-�tB�P~%�T�^���נN6�NV�N�v~� �&f9�D�X� �<AG��C��Z;@�{b�b��p�~�m}K��n~��|���3�!iQ�{�J�Z��:���}���x���NY�s���w���2�Pg�\?�A!�,���j�/�^��,�͟��X��X=�1u��7�u�xӸ�0M_�ER�3�X��V~��*��"*������?�3�i\�M��Ia��� }w
E�O+U~����R`�n�����G%�$ʹ|o�~M�?�"����4�P�K?�"��E�>��x�?a��#!�lZ)�p�?�ρ�Q?B-��\�O��D���������Ǎ�h��S!>aL�����i?�A|&ħ�E|��gC��gB��/��R��ō�"��k �a̅x��A|-�ρ�z�7C�Q%�u��!�_�!�\�� �σ����^�
��a����!~į��� ~-į��Uj�K�7C�-=�o��� �����ײ7�?�0��� ������!~�߫������@�3�⟇�g!�9n��d/�u�a��w �-���oB���.Ŀ����ע����A�W�%��_C�n��^������������C����G ��Z��Q|E?���?ERыb���*�R\�)��>�����\|����t�q2Pq*�R���J�W�D�U�B!T�F+[1L-�˸����`U��'qz��� BI顓@ܒǸ$�&di$�=�Ț�-)(fa�.K�}Yz�e���a�e�K٥Û;��U,�3�h<���x�[�=�en9�o���Y ~�m��n>��r���/�{���@�B�'�/�[�x�c�$��7��� ��ׁ�Z��m���|� ��8�{@���] �	�{A�A!��mmI|;�� �a��# ^�m��O|'�?b�����@� �(����+;�ёz}��bBo:���Л�M?��
�tEi:�2k:ɞ��C���l^yg�n�C�M�z����J��j��
${U�+�U��Zw�3?F�>��{��j����y�����N�7�w���;}��u_�N��v����z�W���ţ3l�Ji-l�s�|�ʎ��,�9�'�yy��M��]㩆&v)�Ig������M��
:�>ܧ�vDL�q��O�V��Mo�n2�m����0'I.ٴ�N8�Ak?YSk#�����;E�J�4Jio�ը�!1r�wD�3%[agZDa�<t�#!�.�mס��֬��%�-�Ԟ��u�[T]�f1h�î�k�kp�+�	����������AQ�LRWT���Y��Í�Ed�V5u�<�kcF���ǜ9zt5���n���t��m={6��1�1�͓1;��<�s���d��R�B���e���B:�WH�ܢ�T?�Ac4�
	n��;IC�R��o{��5���ʎ�4�Ue��e e����;�S��wg�2�tEB����1g�G{������[��5�5�DO!:ky��V�U�MI�<a�<���1�2
3g��ZKa��^��O:|ly'X��A����I�mM��V�>|����0��%9�f>�]|��7�fM�F`�ˬ�-x��}x�]���[6�>5�l`���+x=� �����Ԩ�a���� ���M���-x'��kI�{$E�M�y��d�G1asܒ�wFV��1Z���y�J��g1���{*,q6,q
,q��M_���5fX"�����9�3�>�˒�����@}�^�'�X�s�?ae��9i �B�Й����S�6W�r;ns��K��$޷P�7)7�;$��_$��m�ls���~6i���S
��b|Ix�&Q�_Q������/H0�H�7TX��������Qxn0I�9@��7����D\�m���t�Q��@bp�(nc�O��F���X�ۈD�6��rc,B�7lK⧁�� ~+���
��[��m�B<������B�@�� ~G?�/ �;��]@�|��bK���{��% �
�W��� ~�m�/7��z �X�������
į����F��-��� ��A|3�@|�o���ķ��N��	��w���?į�Q�?Җğ�O�ǃ��@�I ��m�?�|���/���A�� �l.�� �_�ϱ���$�&3��������7؆�k�'�n�ĸ�?� �����@�� �a�U�wْ��A�+ ��<�	Ŀ���6�?c>�o��O �� �#��Ŀ�?���w-B��[�#��	���� ����ۆ��M'�WB�}#H_)e�F���P�|I|�`�7�D����Y��r;�ۜ��&�$�I$�o"��\�MI"�fv!޷���o�gC� ~&���o⧃��A�,?�*�7ؒ�=A�b�;�������E�!~g�_����A�J��W���A|���{Y����lI|�����@�� ��] �`����ķ�xb� >�C ^ �A��%���	�$�$��3�?��������"��+�8ğ�O�'��S@�� �L�E���lI�� �*)���_�/�ۆ��'�'ĸ���o�7���A�m ��E���fK��O��GA�?A� �1��m��|��Ŀ1^�o���@�K ��:�Ŀl�=smI�� �+�)��7����?���O����?���@�/ ���������M�ڑx�8
�O��G������,��M��؅x�0Ӊ�oⷂS(��$�*���'�`~'���J��on�=Q[������s@�?�Ϸ�3�'~�_1�@|%�/�{��� ��W��=�B|�ӮV'~5���׃�:�
�7��F���|��<���x?��@��{@��7��&��dK�� ~-�o�� >j���8�?b��G�����#A�1 �8���VӖz��=�yɩ���I��9�l���`W��cX���J&ڎ��

ￒ$�_B2�/�����\�KI"�e���|����������j@~ ?�_���ϵH�>g�-��������.pu'��\����ެh��f�6��?1��ς��A�� �I���?�K<{N�Y$;&1N)�6�)��r3��av�g�~)j�"�e�U�!�!c��
�i�)��˓��_��e�ɪ�	���h:[#��]F�/XŻ���i�����/l���N�𻌘7��T^�j�~��Hv����'y<m}�ܨyEj͌c��F�C)J�X*k�"�y��M��F��+ݲ��-���,s%�c;�{��HMV�G�cx�,�����e�T�Ͱl�UG%� 
�ވG�-G}w�-;Ɨ�ջꪖT�U�TT��Բ�k�#����bI�iW��d��4�'U���JќsWMA��\�hqpqL�/����s���5� wP�X��#���������;�6��6��̚7��5s��*//�c'?v\�s�n^�wr8�%?��d���Y�Rt����P����3�����/+�ڹ	�,��y	6�];?��P����H�����T�����b1�����U̚�5��_�O|=��97��*�m\��ָ�&�Ԝ��C�q��`;�E}��8b.{���m�����1�?�P�T���&}�� �~nR�~�)��,��y3���	��ӆ.̲]X���0�a����b4�����U��(��Rf�W!�k��}�,;FWՆ9I�ݹ�a���wS�fu�� �ͷ�*��*��*����Ƀ��(U�fZ#��/�m�(�єV/ʬ���er�J�Xe�y�lͶt.ȗRx~I��� ʍLr�I"~P����5�W�E�ؒ[-�K?��&Ǐ���f$�	e�O"Q�	T(~<��oL��I~S*,�Q��2^.���,�?����ߖ���)3~$;��+rj��d�S5�9�)"�AN��bS�Ω[s��ߩ��u��B-������.��z�H���d�G��D6�ذ\W��:~E�W�\��0� �Z�QW�r�����r���.ׅaٜ���pG])���nP�s&mX�V�[�����e~-@>����A���?4�TE����jӕy�5�t��4Ct�R:�HmKva�ݝ&�8�W�]����f���ys���.��f��:���o��W�-'K)b�#����=aM�����Ys�լC_o�/C��>�
E���Z���_Z��!\��$�u���z[�T� 92	/Q���gkk�E��	�b�B\�Ew왣���mml��O�D�Ϻބ[v�(-�Sf-�P�-�mX����eo�Բܠ���%�J�R�,ݰ�a1�`���7�U)�����q1��
�r&I�r
��r2��r:��r*I�r�]NR���~6iy��|
�rĸ�2h��Di��
�r��r	�r)��r9��B�2��%��;@�� �&����j�7��@�����'��?�����B���$��&�Ŀ�_���lC������b|�?������A�� �s��E�oqؒ��@�� �'��G�+����b��g:�C(p�X�ue�:�DiI�jJ�'�ZG��c����,B<��oݒ·N%IZ'����Sn�N��u
IԺ�]�o��|�� �l?���ۃ�Y ~.���gZ�x�-���U ~1���W��2_n��O�
�
b��@|��� ��7���!�ek[��� ��@��{A<g��g�L#>�cC� >��@���A|ć�B�x[,�?�	� �ǀ��@�Ѷ!�0�?ğ1�
���g���A�� �o ��E�矰%��ׁ��@�� �Z5���6�_f>��� Ɲ �����������ۭB���$�9�<�
�?	��O��glC�c���b�������7A�� �]��U��̖���_��/A�7 �? �k������B���$����$�0 ��
�'��A��ۑ���G*��=R)�ͥo�0��Qf�X$;��Rز�G*�)�Zn,7���N���Q���ŰK�Ű�m��Tj?S)�Q$�ܠ3��
� cw����3��/��Le��J.P�I\���*���)'�6;���<����~�R��daN�Z$1h��t�Z��5mla�b)ܻ�X0��݌��Ƥ���̄uH����{���b�jжt�xX�tX�8X���7lK7�6�m����u�D�������eQ��E[lY�eQ�͖E��-��,
ز(`ˢ�-��,
ز(`ˢ�-��,
Vٲ(�ڒxlY�eQ��E[lY~�ٲ(��e1�-�lY`�b [ز��� �,�e1�-��.[�M

�{R00������
]6�(�)�Y ���?��``fq'3
��|XnXn�]��IA壔uQf�0����r�f8���� N/�8�2��L��#�Й�X6g&�T��;UR�mf)p@[��&a�\��e�s�,�
�lK�2�֤�A��4���NШ�7�ѕ�=iҕ�.cx��
����>��1����ѕ��i$k�;xNrɢ9:k�����e��X(t�4E	<K��B��lX��/�"�1h�"�:������Ɔ��/����6,^0AĞ̱a�"#�+=��.l�6p��o��(|p:I܊dN�܂ے\��I��6v��n�~6i�68�w�;P��I���T��<?���D"w���[d����{���A�_�A�R��6ė�O|=�? b�����}A|�_�׀��A|�U����` �A<�A� �[@|�m���'��wB�8�O��� ���@�! ~��Z�x[��
��O�ǃ��@�I ��m�?�|���/���A�� �l.�� �_�ϱ�3mI�M �f����_�o��טO�� ��q?��? ������A�� �^��-�Ŀ�_ �σ��@�� ��lC�3��6��b��?���w@�{ �C�1����Gʇ��k������c�4��k
8�-E	��2~�d�3d�S6�xӚ��Ē��"
�^�mġEN��C(YqX��-/�w5VV��B���V}�K�b�����Hܒ"�S�E$b;��5p e�伻�؇��%��!�����!�2����[�R���9���i�T�w�B��!���eT�2�rYտ�k�mBb9`�(��`E�s˜w��;_��tl�hov�f��Q;�l�ԥ��9�ұUH\�����U�
����S��]b�!�~VTiM��.�����uѡ��}��z�Rz�&l��a��Wr�'lT:�S�'e�k�w�[���%Y�ʬ���ih�/2�+c�|L��9ұ�Y�2��H���^v�e��/7w��U����[������V��|�9\�GW|9[W���m^a��t�LWE*�;�v��E��*e���W��,%�8�UI��8�W����kIҮ�Ј,-mtt�ji�:��{�í��B��+]����.��^�j����9�Z*l����p�����%�e+ip�*ih�(4�����SX����T���؉����ϼ��%�Sf!%j������j&I��'�	5R(fЉ�d<�ka�0,!����qo�%R)��N+�`o V8�0���̱�BF#N+l٫R�����o;���G�C��$��H�Н�[�^�+t7I��.{>B���M��z����OQ�gI���T���$~�I,��z�
z�"��ēlI�{ �}�/��Ŀ�߱�O�g �;���������_��oA�!~�
;�6�·��$m(S��rkDr���DmmC����6��M$1��Sm��(mQ��Ɛ�m�H���I��	Tض�!^\cK⧃� ~k������څ�6�����A�A�. ~'?�� �w��V!~�-���/�KA���_�mC|���7��!ƾ ~��7��� ~? �_e�m�'�-�E��y � ^��>�� �B�� ~�?�GA|�'@|'��Y���d[
�?ğ ��'��A�I�!��?�_1����@�9 �<!��ğk�ŗmI�� �=����	�� �o��ךO�= ����0��������G@�}V!>aK�_��A� �e� �%����Ŀ��1> ���A�� �}���Ŀg�/�%�?���A��@�A�� �{��m���t��)px$�B���(�T�� ?\J�����T��`�?�p;�L��SH��$cx�ޜ�
oF��d�Û�O�� ~�����ۃ�i ~��	�g���!^|ؖ�/�e ~!����	���=lC�.�_�� �
_�k@�^ ~9�_	���{[��mI��{A���@�� �m��7�x�G F�K ��@��� ^�A���%�G���@�a �� �8���m�_g>�'��� �i �L:�?ğ
�� ��X���$�*5���_
���+lC�E�#��b�
�� ���@�- �v'���*�ϱ%�O���A�c �Q�$��?a�6���@�� �k �M�:�Ŀ
�� �o��W�B|�-��
����?�_���A��!�c���K �/ �w�+�����#$��)�x����8���Q}"�X��RD��R��C"C�|y|�O�~�u�LIQ�є�4ɎR�6�'�6��ODI�J-�ODiR�����
�q"Y��^�|"NT}"J\����A�[)z".��uI1\$CT�~�H�v�H���߾�H�v�@��c'5�<.wfB�s�(1A{p��̣�E��f�2�R�V�XY�*�x8IZεs�{�,�_Nbӱ���Ҧ]&J �լ�:L����B�[������k�O�|��ǚ�ʕ�+�j\kj�Xb��H�D��d4WZ`�C�H����(vI��eY�'Ɣ/.B�`�gj���^�;�:���,��T���
U���,C�;6ɐKe�S���wM�(]i%=�`zZ��bR:<�Jwf��H�4�jS�>.���|�o��t\�,=�����K]�#�I?��CQ$\�*��d�5�]͘�뗻�k�$}c���sX�;X�3X�C���2$����x�j�v�
�j�ۮ'slpW�Ū��J���Kޅ�˻�$�$���r�w&��I"y'�L��s��&M��eX�bTQ�2E^B���I|�����r5V����t�-��� �W��U ~?�/�_c���'���ķ�x�s ��[@� �}V!�mK�ׁ�N�1� �kA�!�!��|��'C��@�� �x4�?ğ �O��X��j[��ğ������A��!�o�5��	b\�o �� �׀�����A�� �Z���-��?�������@� �A����?�_�σ���/��g@�s �E���*��iK�?���A�{ �#����6Ŀm>���?B��@�� �� �k�-�������F���P���l�����ߊ��L�9��k�72��DJ)��@J62ب�d3fϖ�H٨��"c�ͦ�2�LB���y#ِ��lmn�ݺ�^jtl�̧H�m��;����avwǺ�[7��Jv�q��}�ܭ�-s6��րi[�T3�ֵƝ�}�U�V�H=`m(`�X[�bV3/a��]��Z�j5GC��rI�&Ɏ���A�h���w����H<KIڷ�1:�Y�ZX����v���j�p�:*`���uV���Ɔ0���u颎N#�[IO�+Ġ�%���y!KIC��G%��wlX��r��ݸ5�^�j��&����-=&!�PRYoJj/�ƨoA:0R�Y5�*a�\����%&^��r{�l�3L�l��զ�u��/�(�{Rf�)��=�������^C��W�������XK�e����un��������^��G����
�~&I�~
��~2��~:��~*I�~�]��OH?����~>n�b\L�_F��_B�j���o��k��Dh��
�~�E�M�����A� �f�����o��כO� �	������?����A�C!��ԖĿ���L/���A�� �5����� ⿀����@��A�� �c�)���d�#/ؒ��@�� �'�#��������3���!�c,��1�2�M�t��Bu%�;��`�H��1T؎aV!�:;߱%��J�tL&;6��:�$W���c�߱���o�@�� ~����@�\?�ϴ����Q	�@�b�'�� �e ��6�/4�� ~���7��:_�kA|=�o�+-B|�[��� ��@��{A<g�]��1�!���m ^�� >
��!>r�-�?���G��c@�Q �h���ğ�υ�g���@�� �L�7�?�*��mI��A�u �*%���_⯱�O�� �>�q'�����o�w���A�� �v�/�w�fu��σ��@�� �Y�4��6�?f>��� �[ ��/�:�Ŀ���oX����$�[���
�	����_ۆ���'�
LbD�At � ��`�!:��f�[�H|t��N$I��I��8�-�	�݈$�nl⣣M'>���1��ۂ���PQ'��
��Ө��--B|h�-�����w�;��]@�N ~g�?�|��A��c	���KA|����@�^ ��"�o^aK� ���}A�j�?�_�����ρ� ��A� �[@��7��V ���ݑ�y�UT*�;�h�۱�1�]K�E�H6n�;�k=���H�Gj�a��a���I}vG2H�$]'SU9������Zυ�yO����$z%E�^e�G��% � q1��4�GEŕn�����y��D��w~I؃N�$�cx�,�����e�T�~X6�?�@M��r���w���<�~4?ʦR�|��E����D����D�����:/)�\�Ӕ��+��r��I����G{7��&��yY�u�L����V!��!��D��,���'
mv�(џ)��H��<�l��N���y�Pv���s��2/{�my�06�"�Ft�0VJQb��56����#����j�����`�
�A�
7�����`�������֔.�)����55�Dv4y�qWc��ES�e9�ۜ9��q͢$���]�N�}x���⃒�z�ES�\���Q���t_$��j����N�^^
	�X���Ey��݇'f�ަ�4#�ڄ]ң~�l�k��GE��|Tl5���K���I�X�[Er�H�X�]�b+��&�G���1bx)���D�qT���ďyH���D�5SacM������K,�ׂ�v�1�⣶!>l>���!�Q �X4���?���GN�:�S^�Y����P{ƅ���P�Dg��I���A������9�o��QòNI�	JW����fy���Ew��L�%ł�^�+�bi�
���0uJC�'���Q�������>v%I��d�]L��.'�b��D��r����lT��P��G��jT�sP��C���@����!;&���SJ����)7sN�2$f���{i#vKq�6b7�����EQb�Pf�;���}\�P�>Iv8U#0���"�$�)6�(�i���G���.|�+�r��r/�r�!�zZ�0����������*��zTv��
ʼ�sR�����F����Q5���xO�3E���#f7���R�;�yg{ŀ��l����H����	\����D!�%�����/fN�c��4'�w��K��cg�<����=�����{�ą�V��T[���6]���A)>8�lU�w����U��#w�4�]�;�,��,�Y7��%�=Y0�_���0��y���e�_?	�o��Y&�������@HȐM�4����J�S�W��T�뻎?��GA����DaB~t69C��9��Wke�B]�M29�2�Fйy�DU���3G̲cp��`��p�S59p}QR�$G�'��^FѪ$�H�86��J<�䈳]�q��oK��Y��!l|;��a�e�I{ ||
�-��&��0�㸣%>�8�OBk�������5"N��#�<e���k�L�S��R����<3M�J�ٛ����G�YU�^�j�<�%�����P�;IV��N�*�S`�歐#P6�2�.fu�ʫ�2��4UQ��T������LU%{JhA4�\!��A�8;�_�0aLf�%M%�ڰ�a�j�j�>.�s�_����]߯�ǎWk�x ҁJ�6�(��\l�[�p]K���&���^�*��tiR-[7�A�]Eqv >ހv�
5��4����q�a�ٴi��To����p���0�&U���w��y�لv��}�1#f�!�(j�6H�˴��Z�&��ݴ���
��?t��Tm�-˨�����p�,9g)o���9#�h���,:����+��d.������(_*o/���j�2��o��W�_h/�m��Y��q�N�䵓F�`Y���󏆪t�,�
QR+��t5������*��HOI�oW���`%P��h+�HZ�&X��F��d�:��
���ɏ��Cr���5l�6⩊*}��vc���l<�1�f���"�@�?�����&.G�iQ�4%�ITV5�(�����/���t�-_�L�ũ����O�?h{��6,'w��XJSǹ�J*��Ԉ�0��V4�L=���襜�L���)�(�mYD�rA��b)���/���4�B�Q�<d�_�s�;kg~43f��y�*��9��� r{��9�oP�5�������T�{H����s�a�9� I��?���^*k�~�*�O�7����_���%��6"i��+f�z�8��ߙ~~<��=�Ԩ�P���JE��|�R��
���
<�}(�"����=/h4�c?�a0Z���VE�b��NN�U{��~����Qͤ��Q��"�sr�PX�F<J�R�I�0R�7V��;+���,��t��q�լq6�Wձ�I��8�V.�t�*[�X5= �TW���5�&L�-?�#���ۭ�X3�T^:=�M�1�sT�V����+#��31�f�x��ߨ3��,K����%�F�p�>g�:4��d�����Aeܢ�U��V���QpV�;k*���L����%ڢi�+kL3���XGŻg;{%S��Zd�ŋ&�]�T������4W�Lja�sZ����i3��ɪWWU����YUW���9���C���t�4C-���8�磌1ws��f:�l�Q�͢�:�xI�G����bX�˨eѼys���|�p*����,��|[�rP����%���4�-�f냱l.��8u��u8��(�7qN��i罜נ�4kK7�h��[���E�TwɬB��p��K��<��Ћ�5���������׋�+<��'��b	�y� *���I3C
>��9��^v˜d�r�k%�x��-D��):3���KCmfwO�I��������V����Ue5�P�䒒�.A�KNcl;�#p�ˣT&��e=�����d�(6��y�; b�!��\�w6��]�,��op�:w�A��&���YUQ����[ۢ}.�y���������f[�2W���`݄\4-k�נFzF�.���3��c�� �Uͼ�G�wOO3�i����-�.+̱LgPt����%��Y��-w@yC�|�L.43?��j�����ԫ�߹zYU]�:�%Z�"��E,�̲�g�R�2�TW.�#7p��:�еoU3MI��--��-�9�7�䢊���Z��X�E���vzy�O)wPV�d�Iʨ�-�%w��r���zkb�@>��65�G�Q�4"�>��$�غp�h m2 ���~l��~F�\l N��RF��_�\}6�tS7%�p|�]i���KT�ƍ��
fCg5%�\�;��>��TCn�iHZ�0�e i��T���&�j�	y+�A��S��s��j��&u���ӆ�O����7�xAV�sbΦ���rz�N�Y�L�����+x����W�s�1���X��;u����i�T�ryy��f)z�"߬qF�v7f�x�4ZB��@�3O!g&��E�-d}+5��g}�s��~I��0oH~.#\_נUq�%�.��tv�v����3�Y�����i�}'�.b׺��L�ݡ��s���� O�Z4-5���*�M|�3֥��������Mힾ�
�|�&~jwK^���>��ۛ���X/��{��@j�Y���^�)R5�ҝ����`jlz0�Z�ܱԄ��TR��R�dX΂æ>��$L���/1X�2�Rc�/0Hv=��`��J��'������	奥BMu=����Sy5S�̛�N�O/�;g>f	����R���˘8��B$�߉��F��''*�	�ǶT>������e���v��v�4k�#c��A��Z�`){���zl?��r��|\��A���������V��s��+���2ƩK��Ӫ��e9�VW7,s���N�[��+e��Z&s�ޙ��Rk$'��M��*]�J=�N}���>,�.uKJ�8� ���{���3��4W�R���|��R��x�����_<#$��/H��.*Z!��E+V�4,��?�XivÜ�wF��k�*�hMUY���FU�����o�1��Ϻ��'΢(��)��_)��ߢ�cRwg$!�6�D+�UO�����:�N��T���d_�BY�Wј|�Y2e`W�TU�j�VTu�����"��R���<ߕg}7B������nU�������¾n�[�U�˺���֭\�U�}�����"(�v���9�U�o,ߧ�kkj���O^�a�J�`�$���;y���}���J��D�`ǯ�u���N��>����-��	���2'���	�)q?�`g��w�T���Ǎ��N���	�W4���H<ʼ���p�ni>ڜP���k��5���>%.GK�<�pZ�+���&��v�<|c>�8)�`���eO]��ƽǦFm�ǰm��2|�ɎA�'ݙ����R�)�W����e��)�)���=����"�b�_v��(���T;���X��M���� ���Y�^?���~�a_)��M��v��)�HceYJ��b�����7w���s³{=��;�ARM����8����璝r��Pmʨ�+iX��{��L5v�؍"��P?Pn�$g�W*a�'�{�a�ו�FO%I�F2�m�LzK�H%L������ם�ƾ�}J|��A\7�"���Gv�օ�|JL�f����FK|��z���WP�Uevm��rTU�\7D���H</(@b�e����R�[ٰBݿ ����A�J�f"�m������&;�j���D$Y$�a�w9�w��Z-;6��*RY���)�h�����R��y�0񉅙����Y�V�+�f1��&{���dW����C/(��������m5Zk{����sS5�1$���ܩS����+�ה��K�nU#��|��u�|��5sLۆ!^ϡe���9�>7|�c�nz�Pz���ş�u�̩�~��mj?1l|_52n9�1�H���e��j�^Po&�m������^zڦtk�Wm�A����$���&qi�H��8)�A��u�{� �Y���U��0�3���2��nz�6t�?l�e��s��oo�f�]��m8���
�F�ױ����lV
�t����w��3����C/̰���aY}
�FB�U������F+���]�M�B�
M��s1eֹ���ܓ�x�u�k[�ɾ����=t-�Pzݬ���J�-/�ν�R�����W�զq(��{ �4��!IK[vI�U�SdGI]-����oH=���ِ��>��%lU4c5�se����ƌgV��9�볉t���ʒ��AJн3K~�\E�2���nR�dN';_�T �&L���i�-��p���r�Vsn�!wc�W��[����5�k/3�(��P���>�)e��}��^�%�M�XH�[S^��d��v��};cJ^�iȫ[%��d4u�հ��r��"�;$6;ٰ������G�<�H�d;t:����G���Wg����Q]�<�}��z�^���ֲ�5]���eu�Ѽ��y"��ȵi�6����|���
jO#s��S͐�]T՞nI����1#�jjU���j*L�۶�
r>
r�����ܘ2u9�UX��F����㆕�����
s
���¨뙽���ZJ9���(�Sf� ه�v`\�v@c��My��������Kf��Y^^�\�|���\�՘�S��oP�η(��7��"S��*����S��F=��bb�I�����|t>:�g�����3����!�t HSGsq ~  t MFUsq ~  t MinorVersionsq ~    t HTRsq ~  t TROsq ~  t DomainIdsq ~    t HTsq ~  t PMajorVersionsq ~     t 
DomainNamet neu_bct HSCLsq ~  t HSCHsq ~  xsr #org.openadaptor.dataobjects.SDOType�s��Ԭ=� Z isPrimitiveJ versionL _uidt Ljava/lang/String;xr 'org.openadaptor.dataobjects.FixedDOTypeDܤ�]ց L _checkedTypesq ~ L 
attributest Ljava/util/Vector;L attributesHashq ~ L nameq ~ :xppsr java.util.Vectorٗ}[�;� I capacityIncrementI elementCount[ elementDatat [Ljava/lang/Object;xp       ur [Ljava.lang.Object;��X�s)l  xp   (sr (org.openadaptor.dataobjects.SDOAttributeJE+���1� L nameq ~ :L typet $Lorg/openadaptor/dataobjects/DOType;xpq ~ sq ~ 9pppt String        q ~ Gsq ~ Cq ~ 
sq ~ 9pppt Int32        q ~ Jsq ~ Cq ~ 'q ~ Isq ~ Cq ~ q ~ Fsq ~ Cq ~ 1q ~ Isq ~ Cq ~ q ~ Isq ~ Cq ~ -q ~ Isq ~ Cq ~ 3q ~ Fsq ~ Cq ~ q ~ Isq ~ Ct Lockedq ~ Fsq ~ Cq ~ q ~ Fsq ~ Cq ~ sq ~ 9pppt Boolean        q ~ Wsq ~ Cq ~ q ~ Vsq ~ Cq ~ q ~ Vsq ~ Cq ~ #q ~ Vsq ~ Cq ~ 5q ~ Vsq ~ Cq ~ 7q ~ Vsq ~ Cq ~ %q ~ Vsq ~ Ct Pswdq ~ Fsq ~ Ct TPq ~ Fsq ~ Cq ~  sq ~ 9pppt Opaque        q ~ dsq ~ Ct CRRulessq ~ 9psq ~ >       uq ~ A   
sq ~ Ct CRKeyq ~ Fsq ~ Ct CRValuesq ~ 9psq ~ >       uq ~ A   
sq ~ Ct Pathq ~ Fsq ~ Ct ANameq ~ Fsq ~ Ct Rulesq ~ 9psq ~ >       uq ~ A   sq ~ Cq ~ vq ~ Fsq ~ Ct Nameq ~ Fsq ~ Ct Descriptionq ~ Fsq ~ Ct AutoGenq ~ Vsq ~ Ct ReadProtq ~ Vsq ~ Ct Whileq ~ Vsq ~ Ct Nocrq ~ Vsq ~ Ct Prtyq ~ Isq ~ Ct InitUseq ~ Isq ~ Ct OnChUseq ~ Vsq ~ Ct OnChOq ~ Vpppppppppxsq ~ ?@     w      q ~ ~q ~ }q ~ vq ~ zq ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ |q ~ {q ~ �q ~ q ~ �q ~ �q ~ �q ~ �xq ~ v         psq ~ Ct SRefq ~ Vsq ~ Ct Aggrq ~ Vsq ~ Ct OrgAttrq ~ Fppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ rq ~ qq ~ tq ~ sq ~ vq ~ uq ~ �q ~ �xt CrossReferenceRule         pppppppppxsq ~ ?@     w      q ~ mq ~ lq ~ kq ~ jxt DomainVersionCrossRefRules         psq ~ Ct OAOsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct OAKq ~ Isq ~ Ct OAVsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct AIDq ~ Fsq ~ Ct AIDAq ~ Fsq ~ Ct ASEq ~ Fsq ~ Ct ASEAq ~ Fppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt OAuthOptions         pppppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �xt DomainVersionOAuthOptions         psq ~ Ct MailInfosq ~ 9psq ~ >       uq ~ A   sq ~ Cq ~ q ~ Fsq ~ Ct INq ~ Fsq ~ Ct MHostq ~ Fsq ~ Ct MUserq ~ Fsq ~ Ct MPswdq ~ Fsq ~ Ct MProtq ~ Isq ~ Ct MPortq ~ Isq ~ Ct MCIq ~ Isq ~ Ct MSSq ~ Vsq ~ Ct SSLq ~ Vsq ~ Ct TLSq ~ Vpppppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt IncomingEmailInfo         psq ~ Ct LINFsq ~ 9psq ~ >       	uq ~ A   
sq ~ Cq ~ q ~ Fsq ~ Ct LCIsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct FLANq ~ Fsq ~ Ct FONq ~ Fsq ~ Ct RFANq ~ Fsq ~ Ct SUONq ~ Fppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt LDAPCorrespondenceInfo         psq ~ Ct AOSLq ~ Vsq ~ Ct CINFq ~ Vsq ~ Ct LATq ~ Isq ~ Ct LFORq ~ Isq ~ Ct FBsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct MPsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct OFq ~ Fsq ~ Ct UAq ~ Fsq ~ Ct PRq ~ Vpppppppxsq ~ ?@     w      q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �xt OAuthMapping         psq ~ Ct UOq ~ Fsq ~ Ct CAq ~ Vpppppppxsq ~ ?@     w      q ~ �q ~ �q ~ q ~ �q ~ �q ~ �xt OAuthLoginOptions         psq ~ Ct GGLq ~ �sq ~ Ct TWq ~ �pxsq ~ ?@     w      	q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~ �q ~q ~q ~ q ~ �q ~ �q ~ �q ~q ~xt 	LoginInfo         psq ~ Ct DBSsq ~ 9psq ~ >       uq ~ A   
sq ~ Cq ~ q ~ Fsq ~ Ct DBq ~ Isq ~ Ct SQLsq ~ 9psq ~ >       uq ~ A   
sq ~ Ct STMTq ~ Fpppppppppxsq ~ ?@     w      q ~q ~xt DatabaseScript_Statement         ppppppppxsq ~ ?@     w      q ~q ~q ~q ~q ~ q ~xt DatabaseScript         psq ~ Cq ~ +q ~ Vsq ~ Cq ~ q ~ Vsq ~ Cq ~ q ~ Vsq ~ Cq ~ /q ~ Vsq ~ Cq ~ )q ~ Vpppppppppxsq ~ ?@     #w   /   q ~ q ~ Yq ~ 
q ~ Hq ~ q ~q ~ �q ~ �q ~ q ~ Xq ~ q ~ Tq ~ q ~ Eq ~
q ~	q ~ q ~ Nq ~ q ~q ~ q ~ Uq ~ q ~ Qq ~ q ~ Lq ~  q ~ bq ~ #q ~ Zq ~ %q ~ ]q ~ 'q ~ Kq ~ )q ~ q ~ +q ~q ~ -q ~ Oq ~ /q ~q ~ �q ~ �q ~ �q ~ �q ~ 1q ~ Mq ~ 3q ~ Pq ~ 5q ~ [q ~ Sq ~ Rq ~ fq ~ eq ~ aq ~ `q ~ 7q ~ \q ~ _q ~ ^xt DomainVersionImpl         p